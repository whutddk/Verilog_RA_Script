/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 7
second: 12
********************************************/

module prm_LUTX1_Po_3_4_4_chk512p2(
	input [2:0] x,
	input [3:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p2
);

	reg [511:0] edge_mask_reg_512p2;
	assign edge_mask_512p2= edge_mask_reg_512p2;

always @( *) begin
    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001101001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001001,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110100011,
11'b11110100100,
11'b11110100101,
11'b11110110100,
11'b11110110101: edge_mask_reg_512p2[0] <= 1'b1;
 		default: edge_mask_reg_512p2[0] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100001,
11'b10010100010: edge_mask_reg_512p2[1] <= 1'b1;
 		default: edge_mask_reg_512p2[1] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100001,
11'b10010100010: edge_mask_reg_512p2[2] <= 1'b1;
 		default: edge_mask_reg_512p2[2] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100001,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110010,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000011,
11'b11011000100,
11'b11110100010,
11'b11110100011,
11'b11110110010,
11'b11110110011,
11'b11110110100,
11'b11111000011,
11'b11111000100: edge_mask_reg_512p2[3] <= 1'b1;
 		default: edge_mask_reg_512p2[3] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[4] <= 1'b1;
 		default: edge_mask_reg_512p2[4] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111001000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b1110111000: edge_mask_reg_512p2[5] <= 1'b1;
 		default: edge_mask_reg_512p2[5] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000010,
11'b11000011,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000010,
11'b111000011,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000: edge_mask_reg_512p2[6] <= 1'b1;
 		default: edge_mask_reg_512p2[6] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110111000,
11'b1110111001,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101: edge_mask_reg_512p2[7] <= 1'b1;
 		default: edge_mask_reg_512p2[7] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100001,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[8] <= 1'b1;
 		default: edge_mask_reg_512p2[8] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[9] <= 1'b1;
 		default: edge_mask_reg_512p2[9] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[10] <= 1'b1;
 		default: edge_mask_reg_512p2[10] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001010011,
11'b10001010100,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b11001110010: edge_mask_reg_512p2[11] <= 1'b1;
 		default: edge_mask_reg_512p2[11] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110100011: edge_mask_reg_512p2[12] <= 1'b1;
 		default: edge_mask_reg_512p2[12] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100: edge_mask_reg_512p2[13] <= 1'b1;
 		default: edge_mask_reg_512p2[13] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100011,
11'b10111100100: edge_mask_reg_512p2[14] <= 1'b1;
 		default: edge_mask_reg_512p2[14] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100: edge_mask_reg_512p2[15] <= 1'b1;
 		default: edge_mask_reg_512p2[15] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111110011,
11'b10111110100: edge_mask_reg_512p2[16] <= 1'b1;
 		default: edge_mask_reg_512p2[16] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010010,
11'b10001010011: edge_mask_reg_512p2[17] <= 1'b1;
 		default: edge_mask_reg_512p2[17] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[18] <= 1'b1;
 		default: edge_mask_reg_512p2[18] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010100011: edge_mask_reg_512p2[19] <= 1'b1;
 		default: edge_mask_reg_512p2[19] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100010101,
11'b1100011000,
11'b1100011001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000010101,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10101000001,
11'b10101000010,
11'b10101000011,
11'b10101000100: edge_mask_reg_512p2[20] <= 1'b1;
 		default: edge_mask_reg_512p2[20] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110011,
11'b10110000100,
11'b10110000101,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110010,
11'b10110110011,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010110011: edge_mask_reg_512p2[21] <= 1'b1;
 		default: edge_mask_reg_512p2[21] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p2[22] <= 1'b1;
 		default: edge_mask_reg_512p2[22] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b10010000000: edge_mask_reg_512p2[23] <= 1'b1;
 		default: edge_mask_reg_512p2[23] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010010000: edge_mask_reg_512p2[24] <= 1'b1;
 		default: edge_mask_reg_512p2[24] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100000,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1100010010,
11'b1100010011,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010011: edge_mask_reg_512p2[25] <= 1'b1;
 		default: edge_mask_reg_512p2[25] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100000,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000100011,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010010,
11'b10001010011: edge_mask_reg_512p2[26] <= 1'b1;
 		default: edge_mask_reg_512p2[26] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100000,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001: edge_mask_reg_512p2[27] <= 1'b1;
 		default: edge_mask_reg_512p2[27] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p2[28] <= 1'b1;
 		default: edge_mask_reg_512p2[28] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p2[29] <= 1'b1;
 		default: edge_mask_reg_512p2[29] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001: edge_mask_reg_512p2[30] <= 1'b1;
 		default: edge_mask_reg_512p2[30] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010: edge_mask_reg_512p2[31] <= 1'b1;
 		default: edge_mask_reg_512p2[31] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[32] <= 1'b1;
 		default: edge_mask_reg_512p2[32] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110010001,
11'b10110010010,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[33] <= 1'b1;
 		default: edge_mask_reg_512p2[33] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[34] <= 1'b1;
 		default: edge_mask_reg_512p2[34] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[35] <= 1'b1;
 		default: edge_mask_reg_512p2[35] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[36] <= 1'b1;
 		default: edge_mask_reg_512p2[36] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[37] <= 1'b1;
 		default: edge_mask_reg_512p2[37] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[38] <= 1'b1;
 		default: edge_mask_reg_512p2[38] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[39] <= 1'b1;
 		default: edge_mask_reg_512p2[39] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[40] <= 1'b1;
 		default: edge_mask_reg_512p2[40] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001011000,
11'b1001011001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b1110100100,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101110010,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011: edge_mask_reg_512p2[41] <= 1'b1;
 		default: edge_mask_reg_512p2[41] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100001,
11'b10010100010,
11'b10101110010,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011: edge_mask_reg_512p2[42] <= 1'b1;
 		default: edge_mask_reg_512p2[42] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100011,
11'b1111100100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100011,
11'b10011100100,
11'b10110110001,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10111000000,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100: edge_mask_reg_512p2[43] <= 1'b1;
 		default: edge_mask_reg_512p2[43] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100100100,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000001,
11'b10101000010,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b11001000010,
11'b11001000011: edge_mask_reg_512p2[44] <= 1'b1;
 		default: edge_mask_reg_512p2[44] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[45] <= 1'b1;
 		default: edge_mask_reg_512p2[45] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[46] <= 1'b1;
 		default: edge_mask_reg_512p2[46] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[47] <= 1'b1;
 		default: edge_mask_reg_512p2[47] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110111000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[48] <= 1'b1;
 		default: edge_mask_reg_512p2[48] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[49] <= 1'b1;
 		default: edge_mask_reg_512p2[49] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[50] <= 1'b1;
 		default: edge_mask_reg_512p2[50] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[51] <= 1'b1;
 		default: edge_mask_reg_512p2[51] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[52] <= 1'b1;
 		default: edge_mask_reg_512p2[52] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p2[53] <= 1'b1;
 		default: edge_mask_reg_512p2[53] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110100,
11'b11010110110,
11'b11010110111,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p2[54] <= 1'b1;
 		default: edge_mask_reg_512p2[54] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11010000111,
11'b11010001000,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p2[55] <= 1'b1;
 		default: edge_mask_reg_512p2[55] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[56] <= 1'b1;
 		default: edge_mask_reg_512p2[56] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[57] <= 1'b1;
 		default: edge_mask_reg_512p2[57] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1011011001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[58] <= 1'b1;
 		default: edge_mask_reg_512p2[58] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[59] <= 1'b1;
 		default: edge_mask_reg_512p2[59] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[60] <= 1'b1;
 		default: edge_mask_reg_512p2[60] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[61] <= 1'b1;
 		default: edge_mask_reg_512p2[61] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[62] <= 1'b1;
 		default: edge_mask_reg_512p2[62] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[63] <= 1'b1;
 		default: edge_mask_reg_512p2[63] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[64] <= 1'b1;
 		default: edge_mask_reg_512p2[64] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[65] <= 1'b1;
 		default: edge_mask_reg_512p2[65] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[66] <= 1'b1;
 		default: edge_mask_reg_512p2[66] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[67] <= 1'b1;
 		default: edge_mask_reg_512p2[67] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[68] <= 1'b1;
 		default: edge_mask_reg_512p2[68] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[69] <= 1'b1;
 		default: edge_mask_reg_512p2[69] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[70] <= 1'b1;
 		default: edge_mask_reg_512p2[70] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[71] <= 1'b1;
 		default: edge_mask_reg_512p2[71] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[72] <= 1'b1;
 		default: edge_mask_reg_512p2[72] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[73] <= 1'b1;
 		default: edge_mask_reg_512p2[73] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[74] <= 1'b1;
 		default: edge_mask_reg_512p2[74] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[75] <= 1'b1;
 		default: edge_mask_reg_512p2[75] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[76] <= 1'b1;
 		default: edge_mask_reg_512p2[76] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[77] <= 1'b1;
 		default: edge_mask_reg_512p2[77] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001011000,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[78] <= 1'b1;
 		default: edge_mask_reg_512p2[78] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[79] <= 1'b1;
 		default: edge_mask_reg_512p2[79] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010010,
11'b1010011,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[80] <= 1'b1;
 		default: edge_mask_reg_512p2[80] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010010,
11'b1010011,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010010,
11'b1001010011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[81] <= 1'b1;
 		default: edge_mask_reg_512p2[81] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010010,
11'b1010011,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[82] <= 1'b1;
 		default: edge_mask_reg_512p2[82] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110000011,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100001,
11'b10110100010,
11'b10110110001,
11'b10110110010: edge_mask_reg_512p2[83] <= 1'b1;
 		default: edge_mask_reg_512p2[83] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100011000,
11'b1100011001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11100000011,
11'b11100000100: edge_mask_reg_512p2[84] <= 1'b1;
 		default: edge_mask_reg_512p2[84] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100011000,
11'b1100011001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11100000011,
11'b11100000100: edge_mask_reg_512p2[85] <= 1'b1;
 		default: edge_mask_reg_512p2[85] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1100000100,
11'b1100000101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10100000000,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b11000000001,
11'b11000000010,
11'b11000000011,
11'b11000000100: edge_mask_reg_512p2[86] <= 1'b1;
 		default: edge_mask_reg_512p2[86] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100011000,
11'b1100011001,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100110001,
11'b10101000001: edge_mask_reg_512p2[87] <= 1'b1;
 		default: edge_mask_reg_512p2[87] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010011,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[88] <= 1'b1;
 		default: edge_mask_reg_512p2[88] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010011,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[89] <= 1'b1;
 		default: edge_mask_reg_512p2[89] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010010,
11'b1111010011,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[90] <= 1'b1;
 		default: edge_mask_reg_512p2[90] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011010010,
11'b10011010011: edge_mask_reg_512p2[91] <= 1'b1;
 		default: edge_mask_reg_512p2[91] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011010010,
11'b10011010011,
11'b10011010100: edge_mask_reg_512p2[92] <= 1'b1;
 		default: edge_mask_reg_512p2[92] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111101000,
11'b1111101001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011010010,
11'b10011010011,
11'b10011010100: edge_mask_reg_512p2[93] <= 1'b1;
 		default: edge_mask_reg_512p2[93] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111101000,
11'b1111101001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101: edge_mask_reg_512p2[94] <= 1'b1;
 		default: edge_mask_reg_512p2[94] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111101000,
11'b1111101001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100010,
11'b10011100011,
11'b10011100100: edge_mask_reg_512p2[95] <= 1'b1;
 		default: edge_mask_reg_512p2[95] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[96] <= 1'b1;
 		default: edge_mask_reg_512p2[96] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p2[97] <= 1'b1;
 		default: edge_mask_reg_512p2[97] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[98] <= 1'b1;
 		default: edge_mask_reg_512p2[98] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110010001: edge_mask_reg_512p2[99] <= 1'b1;
 		default: edge_mask_reg_512p2[99] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011: edge_mask_reg_512p2[100] <= 1'b1;
 		default: edge_mask_reg_512p2[100] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[101] <= 1'b1;
 		default: edge_mask_reg_512p2[101] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[102] <= 1'b1;
 		default: edge_mask_reg_512p2[102] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[103] <= 1'b1;
 		default: edge_mask_reg_512p2[103] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[104] <= 1'b1;
 		default: edge_mask_reg_512p2[104] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010000,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100111,
11'b1111101000,
11'b10010110001,
11'b10010110010,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011010001,
11'b10011010010,
11'b10011010011: edge_mask_reg_512p2[105] <= 1'b1;
 		default: edge_mask_reg_512p2[105] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100011000,
11'b1100011001,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000001000,
11'b10000010110,
11'b10000010111,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11100000011,
11'b11100000100,
11'b11100000101: edge_mask_reg_512p2[106] <= 1'b1;
 		default: edge_mask_reg_512p2[106] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000: edge_mask_reg_512p2[107] <= 1'b1;
 		default: edge_mask_reg_512p2[107] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110011: edge_mask_reg_512p2[108] <= 1'b1;
 		default: edge_mask_reg_512p2[108] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010011: edge_mask_reg_512p2[109] <= 1'b1;
 		default: edge_mask_reg_512p2[109] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[110] <= 1'b1;
 		default: edge_mask_reg_512p2[110] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p2[111] <= 1'b1;
 		default: edge_mask_reg_512p2[111] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p2[112] <= 1'b1;
 		default: edge_mask_reg_512p2[112] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101010000,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p2[113] <= 1'b1;
 		default: edge_mask_reg_512p2[113] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11000110,
11'b11000111,
11'b11001000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10011110110,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111110000,
11'b10111110001,
11'b10111110010,
11'b10111110011,
11'b10111110100,
11'b10111110101,
11'b11011110000,
11'b11011110001,
11'b11011110010,
11'b11011110011: edge_mask_reg_512p2[114] <= 1'b1;
 		default: edge_mask_reg_512p2[114] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11101010010,
11'b11101010011,
11'b11101100010,
11'b11101100011,
11'b11101100100,
11'b11101110010,
11'b11101110011: edge_mask_reg_512p2[115] <= 1'b1;
 		default: edge_mask_reg_512p2[115] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101100110,
11'b1101100111,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010010,
11'b10110010011,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101: edge_mask_reg_512p2[116] <= 1'b1;
 		default: edge_mask_reg_512p2[116] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010110111,
11'b1010111000,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110000,
11'b1111110001,
11'b1111110010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111110000,
11'b10111110001,
11'b10111110010,
11'b10111110011: edge_mask_reg_512p2[117] <= 1'b1;
 		default: edge_mask_reg_512p2[117] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110: edge_mask_reg_512p2[118] <= 1'b1;
 		default: edge_mask_reg_512p2[118] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101000,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000011,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11101010011,
11'b11101010100,
11'b11101010101,
11'b11101100011,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[119] <= 1'b1;
 		default: edge_mask_reg_512p2[119] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p2[120] <= 1'b1;
 		default: edge_mask_reg_512p2[120] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p2[121] <= 1'b1;
 		default: edge_mask_reg_512p2[121] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100010: edge_mask_reg_512p2[122] <= 1'b1;
 		default: edge_mask_reg_512p2[122] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100010: edge_mask_reg_512p2[123] <= 1'b1;
 		default: edge_mask_reg_512p2[123] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100010: edge_mask_reg_512p2[124] <= 1'b1;
 		default: edge_mask_reg_512p2[124] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[125] <= 1'b1;
 		default: edge_mask_reg_512p2[125] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[126] <= 1'b1;
 		default: edge_mask_reg_512p2[126] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[127] <= 1'b1;
 		default: edge_mask_reg_512p2[127] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010,
11'b10110100010: edge_mask_reg_512p2[128] <= 1'b1;
 		default: edge_mask_reg_512p2[128] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100010,
11'b10010100011: edge_mask_reg_512p2[129] <= 1'b1;
 		default: edge_mask_reg_512p2[129] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100010,
11'b10010100011: edge_mask_reg_512p2[130] <= 1'b1;
 		default: edge_mask_reg_512p2[130] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100010,
11'b10010100011: edge_mask_reg_512p2[131] <= 1'b1;
 		default: edge_mask_reg_512p2[131] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110100,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111001,
11'b10001110100,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10110010100: edge_mask_reg_512p2[132] <= 1'b1;
 		default: edge_mask_reg_512p2[132] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110010,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000011,
11'b11011000100,
11'b11110010011,
11'b11110010100,
11'b11110100011,
11'b11110100100,
11'b11110110011,
11'b11110110100,
11'b11111000011,
11'b11111000100: edge_mask_reg_512p2[133] <= 1'b1;
 		default: edge_mask_reg_512p2[133] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[134] <= 1'b1;
 		default: edge_mask_reg_512p2[134] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b1110011001,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000011,
11'b10010000100: edge_mask_reg_512p2[135] <= 1'b1;
 		default: edge_mask_reg_512p2[135] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100010101,
11'b1100011000,
11'b1100011001,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000010101,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000001,
11'b10101000010,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b11000110010,
11'b11000110011,
11'b11001000010,
11'b11001000011: edge_mask_reg_512p2[136] <= 1'b1;
 		default: edge_mask_reg_512p2[136] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[137] <= 1'b1;
 		default: edge_mask_reg_512p2[137] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[138] <= 1'b1;
 		default: edge_mask_reg_512p2[138] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[139] <= 1'b1;
 		default: edge_mask_reg_512p2[139] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[140] <= 1'b1;
 		default: edge_mask_reg_512p2[140] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[141] <= 1'b1;
 		default: edge_mask_reg_512p2[141] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[142] <= 1'b1;
 		default: edge_mask_reg_512p2[142] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[143] <= 1'b1;
 		default: edge_mask_reg_512p2[143] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[144] <= 1'b1;
 		default: edge_mask_reg_512p2[144] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[145] <= 1'b1;
 		default: edge_mask_reg_512p2[145] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[146] <= 1'b1;
 		default: edge_mask_reg_512p2[146] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[147] <= 1'b1;
 		default: edge_mask_reg_512p2[147] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[148] <= 1'b1;
 		default: edge_mask_reg_512p2[148] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[149] <= 1'b1;
 		default: edge_mask_reg_512p2[149] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[150] <= 1'b1;
 		default: edge_mask_reg_512p2[150] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[151] <= 1'b1;
 		default: edge_mask_reg_512p2[151] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[152] <= 1'b1;
 		default: edge_mask_reg_512p2[152] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[153] <= 1'b1;
 		default: edge_mask_reg_512p2[153] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[154] <= 1'b1;
 		default: edge_mask_reg_512p2[154] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[155] <= 1'b1;
 		default: edge_mask_reg_512p2[155] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[156] <= 1'b1;
 		default: edge_mask_reg_512p2[156] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[157] <= 1'b1;
 		default: edge_mask_reg_512p2[157] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[158] <= 1'b1;
 		default: edge_mask_reg_512p2[158] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[159] <= 1'b1;
 		default: edge_mask_reg_512p2[159] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[160] <= 1'b1;
 		default: edge_mask_reg_512p2[160] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[161] <= 1'b1;
 		default: edge_mask_reg_512p2[161] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[162] <= 1'b1;
 		default: edge_mask_reg_512p2[162] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[163] <= 1'b1;
 		default: edge_mask_reg_512p2[163] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100010,
11'b1001100011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[164] <= 1'b1;
 		default: edge_mask_reg_512p2[164] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100010,
11'b1001100011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[165] <= 1'b1;
 		default: edge_mask_reg_512p2[165] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111001000,
11'b1001100010,
11'b1001100011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011001000,
11'b1011001001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[166] <= 1'b1;
 		default: edge_mask_reg_512p2[166] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[167] <= 1'b1;
 		default: edge_mask_reg_512p2[167] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110010010,
11'b10110010011,
11'b10110100011: edge_mask_reg_512p2[168] <= 1'b1;
 		default: edge_mask_reg_512p2[168] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101000,
11'b1100101001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000010010,
11'b11000010011,
11'b11000010100,
11'b11000010101,
11'b11100000010,
11'b11100000011: edge_mask_reg_512p2[169] <= 1'b1;
 		default: edge_mask_reg_512p2[169] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101000,
11'b1100101001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000010010,
11'b11000010011,
11'b11000010100,
11'b11000010101,
11'b11100000010,
11'b11100000011: edge_mask_reg_512p2[170] <= 1'b1;
 		default: edge_mask_reg_512p2[170] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101000,
11'b1100101001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000001000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11000010010,
11'b11000010011,
11'b11000010100,
11'b11000010101,
11'b11100000010,
11'b11100000011,
11'b11100000100: edge_mask_reg_512p2[171] <= 1'b1;
 		default: edge_mask_reg_512p2[171] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101000,
11'b1100101001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000001000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010010,
11'b11000010011,
11'b11000010100,
11'b11000010101,
11'b11000010110,
11'b11100000010,
11'b11100000011,
11'b11100000100,
11'b11100000101: edge_mask_reg_512p2[172] <= 1'b1;
 		default: edge_mask_reg_512p2[172] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[173] <= 1'b1;
 		default: edge_mask_reg_512p2[173] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[174] <= 1'b1;
 		default: edge_mask_reg_512p2[174] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010010: edge_mask_reg_512p2[175] <= 1'b1;
 		default: edge_mask_reg_512p2[175] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[176] <= 1'b1;
 		default: edge_mask_reg_512p2[176] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[177] <= 1'b1;
 		default: edge_mask_reg_512p2[177] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[178] <= 1'b1;
 		default: edge_mask_reg_512p2[178] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[179] <= 1'b1;
 		default: edge_mask_reg_512p2[179] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[180] <= 1'b1;
 		default: edge_mask_reg_512p2[180] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101000011,
11'b10101000100,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100010,
11'b11001110010: edge_mask_reg_512p2[181] <= 1'b1;
 		default: edge_mask_reg_512p2[181] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000011,
11'b10101000100,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[182] <= 1'b1;
 		default: edge_mask_reg_512p2[182] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[183] <= 1'b1;
 		default: edge_mask_reg_512p2[183] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[184] <= 1'b1;
 		default: edge_mask_reg_512p2[184] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[185] <= 1'b1;
 		default: edge_mask_reg_512p2[185] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[186] <= 1'b1;
 		default: edge_mask_reg_512p2[186] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[187] <= 1'b1;
 		default: edge_mask_reg_512p2[187] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11101110011: edge_mask_reg_512p2[188] <= 1'b1;
 		default: edge_mask_reg_512p2[188] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010100,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11101110010,
11'b11101110011: edge_mask_reg_512p2[189] <= 1'b1;
 		default: edge_mask_reg_512p2[189] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11101110011: edge_mask_reg_512p2[190] <= 1'b1;
 		default: edge_mask_reg_512p2[190] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110: edge_mask_reg_512p2[191] <= 1'b1;
 		default: edge_mask_reg_512p2[191] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11101100011,
11'b11101100100: edge_mask_reg_512p2[192] <= 1'b1;
 		default: edge_mask_reg_512p2[192] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110101000,
11'b1110101001,
11'b10010000001: edge_mask_reg_512p2[193] <= 1'b1;
 		default: edge_mask_reg_512p2[193] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010110011,
11'b11010110100: edge_mask_reg_512p2[194] <= 1'b1;
 		default: edge_mask_reg_512p2[194] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[195] <= 1'b1;
 		default: edge_mask_reg_512p2[195] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[196] <= 1'b1;
 		default: edge_mask_reg_512p2[196] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[197] <= 1'b1;
 		default: edge_mask_reg_512p2[197] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b10010000000,
11'b10010000001,
11'b10010010000: edge_mask_reg_512p2[198] <= 1'b1;
 		default: edge_mask_reg_512p2[198] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[199] <= 1'b1;
 		default: edge_mask_reg_512p2[199] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[200] <= 1'b1;
 		default: edge_mask_reg_512p2[200] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[201] <= 1'b1;
 		default: edge_mask_reg_512p2[201] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[202] <= 1'b1;
 		default: edge_mask_reg_512p2[202] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[203] <= 1'b1;
 		default: edge_mask_reg_512p2[203] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110001000,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010001000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[204] <= 1'b1;
 		default: edge_mask_reg_512p2[204] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[205] <= 1'b1;
 		default: edge_mask_reg_512p2[205] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101111000,
11'b10001000010,
11'b10001000011,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011: edge_mask_reg_512p2[206] <= 1'b1;
 		default: edge_mask_reg_512p2[206] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011: edge_mask_reg_512p2[207] <= 1'b1;
 		default: edge_mask_reg_512p2[207] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100010,
11'b10001100011: edge_mask_reg_512p2[208] <= 1'b1;
 		default: edge_mask_reg_512p2[208] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110010,
11'b10000110011,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100010,
11'b10001100011: edge_mask_reg_512p2[209] <= 1'b1;
 		default: edge_mask_reg_512p2[209] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[210] <= 1'b1;
 		default: edge_mask_reg_512p2[210] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1100100100,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010011: edge_mask_reg_512p2[211] <= 1'b1;
 		default: edge_mask_reg_512p2[211] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000011011,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b11000010010,
11'b11000010011: edge_mask_reg_512p2[212] <= 1'b1;
 		default: edge_mask_reg_512p2[212] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11101010100,
11'b11101100011,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[213] <= 1'b1;
 		default: edge_mask_reg_512p2[213] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11101010011,
11'b11101010100,
11'b11101100011,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[214] <= 1'b1;
 		default: edge_mask_reg_512p2[214] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000: edge_mask_reg_512p2[215] <= 1'b1;
 		default: edge_mask_reg_512p2[215] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[216] <= 1'b1;
 		default: edge_mask_reg_512p2[216] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110001,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11101010010,
11'b11101010011,
11'b11101100010,
11'b11101100011,
11'b11101100100,
11'b11101110010,
11'b11101110011: edge_mask_reg_512p2[217] <= 1'b1;
 		default: edge_mask_reg_512p2[217] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001001,
11'b110001010,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100100,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p2[218] <= 1'b1;
 		default: edge_mask_reg_512p2[218] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[219] <= 1'b1;
 		default: edge_mask_reg_512p2[219] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101110010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[220] <= 1'b1;
 		default: edge_mask_reg_512p2[220] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011: edge_mask_reg_512p2[221] <= 1'b1;
 		default: edge_mask_reg_512p2[221] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010010011,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[222] <= 1'b1;
 		default: edge_mask_reg_512p2[222] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p2[223] <= 1'b1;
 		default: edge_mask_reg_512p2[223] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p2[224] <= 1'b1;
 		default: edge_mask_reg_512p2[224] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p2[225] <= 1'b1;
 		default: edge_mask_reg_512p2[225] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111001000,
11'b1111001001,
11'b1111010010,
11'b1111010011,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[226] <= 1'b1;
 		default: edge_mask_reg_512p2[226] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10110100001: edge_mask_reg_512p2[227] <= 1'b1;
 		default: edge_mask_reg_512p2[227] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100: edge_mask_reg_512p2[228] <= 1'b1;
 		default: edge_mask_reg_512p2[228] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100101000,
11'b1100101001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[229] <= 1'b1;
 		default: edge_mask_reg_512p2[229] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010001000,
11'b1010001001,
11'b1100101000,
11'b1100101001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[230] <= 1'b1;
 		default: edge_mask_reg_512p2[230] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p2[231] <= 1'b1;
 		default: edge_mask_reg_512p2[231] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10101100,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b10111100,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11001011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010110011,
11'b11010110100: edge_mask_reg_512p2[232] <= 1'b1;
 		default: edge_mask_reg_512p2[232] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110011,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110001,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010100001,
11'b11010100010,
11'b11010100011,
11'b11010110001,
11'b11010110010: edge_mask_reg_512p2[233] <= 1'b1;
 		default: edge_mask_reg_512p2[233] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110011,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110001,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100001,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010110001,
11'b11010110010: edge_mask_reg_512p2[234] <= 1'b1;
 		default: edge_mask_reg_512p2[234] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p2[235] <= 1'b1;
 		default: edge_mask_reg_512p2[235] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10111000,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10101110011,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110010001: edge_mask_reg_512p2[236] <= 1'b1;
 		default: edge_mask_reg_512p2[236] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[237] <= 1'b1;
 		default: edge_mask_reg_512p2[237] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[238] <= 1'b1;
 		default: edge_mask_reg_512p2[238] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[239] <= 1'b1;
 		default: edge_mask_reg_512p2[239] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p2[240] <= 1'b1;
 		default: edge_mask_reg_512p2[240] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111011000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p2[241] <= 1'b1;
 		default: edge_mask_reg_512p2[241] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11110100011,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p2[242] <= 1'b1;
 		default: edge_mask_reg_512p2[242] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p2[243] <= 1'b1;
 		default: edge_mask_reg_512p2[243] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11110010011,
11'b11110010100,
11'b11110010101,
11'b11110100011,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p2[244] <= 1'b1;
 		default: edge_mask_reg_512p2[244] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p2[245] <= 1'b1;
 		default: edge_mask_reg_512p2[245] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10110010001: edge_mask_reg_512p2[246] <= 1'b1;
 		default: edge_mask_reg_512p2[246] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[247] <= 1'b1;
 		default: edge_mask_reg_512p2[247] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[248] <= 1'b1;
 		default: edge_mask_reg_512p2[248] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110111000,
11'b1110111001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010: edge_mask_reg_512p2[249] <= 1'b1;
 		default: edge_mask_reg_512p2[249] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110110,
11'b1101110111,
11'b1101111001,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001000101,
11'b11001000110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110: edge_mask_reg_512p2[250] <= 1'b1;
 		default: edge_mask_reg_512p2[250] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010: edge_mask_reg_512p2[251] <= 1'b1;
 		default: edge_mask_reg_512p2[251] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[252] <= 1'b1;
 		default: edge_mask_reg_512p2[252] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[253] <= 1'b1;
 		default: edge_mask_reg_512p2[253] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101: edge_mask_reg_512p2[254] <= 1'b1;
 		default: edge_mask_reg_512p2[254] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010110111,
11'b1010111000,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110000,
11'b1111110001,
11'b1111110010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111110010,
11'b10111110011: edge_mask_reg_512p2[255] <= 1'b1;
 		default: edge_mask_reg_512p2[255] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b1110101001,
11'b10001100101,
11'b10001100110,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101: edge_mask_reg_512p2[256] <= 1'b1;
 		default: edge_mask_reg_512p2[256] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110101: edge_mask_reg_512p2[257] <= 1'b1;
 		default: edge_mask_reg_512p2[257] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[258] <= 1'b1;
 		default: edge_mask_reg_512p2[258] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[259] <= 1'b1;
 		default: edge_mask_reg_512p2[259] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[260] <= 1'b1;
 		default: edge_mask_reg_512p2[260] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010101,
11'b11001010110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11110000011: edge_mask_reg_512p2[261] <= 1'b1;
 		default: edge_mask_reg_512p2[261] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010001,
11'b10010010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b10010000000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000: edge_mask_reg_512p2[262] <= 1'b1;
 		default: edge_mask_reg_512p2[262] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1101110010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110111,
11'b1110111000: edge_mask_reg_512p2[263] <= 1'b1;
 		default: edge_mask_reg_512p2[263] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11001011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000111,
11'b10111001000,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000111,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110100111,
11'b11110110100,
11'b11110110101,
11'b11110110110,
11'b11110110111,
11'b11110111000,
11'b11111000101: edge_mask_reg_512p2[264] <= 1'b1;
 		default: edge_mask_reg_512p2[264] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100011,
11'b10110100100,
11'b10110110000,
11'b10110110001,
11'b10110110011,
11'b10110110100,
11'b10111000001: edge_mask_reg_512p2[265] <= 1'b1;
 		default: edge_mask_reg_512p2[265] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000: edge_mask_reg_512p2[266] <= 1'b1;
 		default: edge_mask_reg_512p2[266] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[267] <= 1'b1;
 		default: edge_mask_reg_512p2[267] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000101,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[268] <= 1'b1;
 		default: edge_mask_reg_512p2[268] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[269] <= 1'b1;
 		default: edge_mask_reg_512p2[269] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[270] <= 1'b1;
 		default: edge_mask_reg_512p2[270] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010111,
11'b111011000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100011: edge_mask_reg_512p2[271] <= 1'b1;
 		default: edge_mask_reg_512p2[271] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[272] <= 1'b1;
 		default: edge_mask_reg_512p2[272] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[273] <= 1'b1;
 		default: edge_mask_reg_512p2[273] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[274] <= 1'b1;
 		default: edge_mask_reg_512p2[274] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[275] <= 1'b1;
 		default: edge_mask_reg_512p2[275] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[276] <= 1'b1;
 		default: edge_mask_reg_512p2[276] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[277] <= 1'b1;
 		default: edge_mask_reg_512p2[277] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[278] <= 1'b1;
 		default: edge_mask_reg_512p2[278] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[279] <= 1'b1;
 		default: edge_mask_reg_512p2[279] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[280] <= 1'b1;
 		default: edge_mask_reg_512p2[280] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010100001,
11'b10010110001: edge_mask_reg_512p2[281] <= 1'b1;
 		default: edge_mask_reg_512p2[281] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110100010,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p2[282] <= 1'b1;
 		default: edge_mask_reg_512p2[282] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000100,
11'b1001000101,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001011000,
11'b1001011001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101001000,
11'b1101001001,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[283] <= 1'b1;
 		default: edge_mask_reg_512p2[283] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001011000,
11'b1001011001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101001000,
11'b1101001001,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[284] <= 1'b1;
 		default: edge_mask_reg_512p2[284] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101001000,
11'b1101001001,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[285] <= 1'b1;
 		default: edge_mask_reg_512p2[285] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000100,
11'b1100000101,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b10000000100,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[286] <= 1'b1;
 		default: edge_mask_reg_512p2[286] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000100,
11'b1100000101,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000011,
11'b10100000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[287] <= 1'b1;
 		default: edge_mask_reg_512p2[287] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000011,
11'b10100000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[288] <= 1'b1;
 		default: edge_mask_reg_512p2[288] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[289] <= 1'b1;
 		default: edge_mask_reg_512p2[289] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[290] <= 1'b1;
 		default: edge_mask_reg_512p2[290] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b11000000010,
11'b11000010010: edge_mask_reg_512p2[291] <= 1'b1;
 		default: edge_mask_reg_512p2[291] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110110001: edge_mask_reg_512p2[292] <= 1'b1;
 		default: edge_mask_reg_512p2[292] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1101000,
11'b1101001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101001001,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b11000100010,
11'b11000110010,
11'b11000110011: edge_mask_reg_512p2[293] <= 1'b1;
 		default: edge_mask_reg_512p2[293] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100001,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010110010,
11'b11010110011: edge_mask_reg_512p2[294] <= 1'b1;
 		default: edge_mask_reg_512p2[294] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[295] <= 1'b1;
 		default: edge_mask_reg_512p2[295] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[296] <= 1'b1;
 		default: edge_mask_reg_512p2[296] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1011011001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[297] <= 1'b1;
 		default: edge_mask_reg_512p2[297] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[298] <= 1'b1;
 		default: edge_mask_reg_512p2[298] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b1110110011,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[299] <= 1'b1;
 		default: edge_mask_reg_512p2[299] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10101110001,
11'b10110000001: edge_mask_reg_512p2[300] <= 1'b1;
 		default: edge_mask_reg_512p2[300] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10110100010,
11'b10110100011,
11'b10110110000,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10111000000,
11'b10111000001: edge_mask_reg_512p2[301] <= 1'b1;
 		default: edge_mask_reg_512p2[301] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010010000,
11'b10010010001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[302] <= 1'b1;
 		default: edge_mask_reg_512p2[302] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[303] <= 1'b1;
 		default: edge_mask_reg_512p2[303] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[304] <= 1'b1;
 		default: edge_mask_reg_512p2[304] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000010,
11'b1011000011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[305] <= 1'b1;
 		default: edge_mask_reg_512p2[305] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[306] <= 1'b1;
 		default: edge_mask_reg_512p2[306] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[307] <= 1'b1;
 		default: edge_mask_reg_512p2[307] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[308] <= 1'b1;
 		default: edge_mask_reg_512p2[308] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[309] <= 1'b1;
 		default: edge_mask_reg_512p2[309] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111001000,
11'b1111001001,
11'b10010010011,
11'b10010010100,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[310] <= 1'b1;
 		default: edge_mask_reg_512p2[310] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001,
11'b10010010001,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[311] <= 1'b1;
 		default: edge_mask_reg_512p2[311] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101000011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101011000,
11'b1101011001,
11'b1101101000,
11'b1101101001,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[312] <= 1'b1;
 		default: edge_mask_reg_512p2[312] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001010011,
11'b10001010100,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011,
11'b11010000010: edge_mask_reg_512p2[313] <= 1'b1;
 		default: edge_mask_reg_512p2[313] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001110010,
11'b11001110011,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p2[314] <= 1'b1;
 		default: edge_mask_reg_512p2[314] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001110010,
11'b11010000010: edge_mask_reg_512p2[315] <= 1'b1;
 		default: edge_mask_reg_512p2[315] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011001,
11'b1011011010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111001,
11'b1110111010,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110100010,
11'b10110100011,
11'b10110110010,
11'b10110110011: edge_mask_reg_512p2[316] <= 1'b1;
 		default: edge_mask_reg_512p2[316] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101: edge_mask_reg_512p2[317] <= 1'b1;
 		default: edge_mask_reg_512p2[317] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p2[318] <= 1'b1;
 		default: edge_mask_reg_512p2[318] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10110100001: edge_mask_reg_512p2[319] <= 1'b1;
 		default: edge_mask_reg_512p2[319] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001111000,
11'b1001111001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[320] <= 1'b1;
 		default: edge_mask_reg_512p2[320] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110000010,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110100,
11'b1110111000,
11'b1110111001,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[321] <= 1'b1;
 		default: edge_mask_reg_512p2[321] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000011,
11'b11011000100,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11110100011,
11'b11110100100,
11'b11110100101,
11'b11110110011,
11'b11110110100,
11'b11110110101,
11'b11111000011: edge_mask_reg_512p2[322] <= 1'b1;
 		default: edge_mask_reg_512p2[322] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p2[323] <= 1'b1;
 		default: edge_mask_reg_512p2[323] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[324] <= 1'b1;
 		default: edge_mask_reg_512p2[324] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[325] <= 1'b1;
 		default: edge_mask_reg_512p2[325] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110000000,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100011: edge_mask_reg_512p2[326] <= 1'b1;
 		default: edge_mask_reg_512p2[326] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110000000,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100: edge_mask_reg_512p2[327] <= 1'b1;
 		default: edge_mask_reg_512p2[327] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010000,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[328] <= 1'b1;
 		default: edge_mask_reg_512p2[328] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001001,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101001000,
11'b1101001001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100: edge_mask_reg_512p2[329] <= 1'b1;
 		default: edge_mask_reg_512p2[329] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001001,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100110011,
11'b10100110100: edge_mask_reg_512p2[330] <= 1'b1;
 		default: edge_mask_reg_512p2[330] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101001000,
11'b101001001,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001001,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101: edge_mask_reg_512p2[331] <= 1'b1;
 		default: edge_mask_reg_512p2[331] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001001,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101: edge_mask_reg_512p2[332] <= 1'b1;
 		default: edge_mask_reg_512p2[332] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11001000,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11110010011,
11'b11110010100: edge_mask_reg_512p2[333] <= 1'b1;
 		default: edge_mask_reg_512p2[333] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101: edge_mask_reg_512p2[334] <= 1'b1;
 		default: edge_mask_reg_512p2[334] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001001,
11'b110001010,
11'b1000101000,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001001,
11'b1010001010,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101100111: edge_mask_reg_512p2[335] <= 1'b1;
 		default: edge_mask_reg_512p2[335] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110001,
11'b10010110010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101: edge_mask_reg_512p2[336] <= 1'b1;
 		default: edge_mask_reg_512p2[336] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11001000100,
11'b11001000101,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11101010010,
11'b11101010011,
11'b11101010100,
11'b11101100010,
11'b11101100011,
11'b11101100100: edge_mask_reg_512p2[337] <= 1'b1;
 		default: edge_mask_reg_512p2[337] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110100111,
11'b110101000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110010,
11'b10111110011,
11'b11011010011,
11'b11011010100: edge_mask_reg_512p2[338] <= 1'b1;
 		default: edge_mask_reg_512p2[338] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010: edge_mask_reg_512p2[339] <= 1'b1;
 		default: edge_mask_reg_512p2[339] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p2[340] <= 1'b1;
 		default: edge_mask_reg_512p2[340] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p2[341] <= 1'b1;
 		default: edge_mask_reg_512p2[341] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p2[342] <= 1'b1;
 		default: edge_mask_reg_512p2[342] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10111000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101: edge_mask_reg_512p2[343] <= 1'b1;
 		default: edge_mask_reg_512p2[343] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001001000,
11'b1001001001,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010101: edge_mask_reg_512p2[344] <= 1'b1;
 		default: edge_mask_reg_512p2[344] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101: edge_mask_reg_512p2[345] <= 1'b1;
 		default: edge_mask_reg_512p2[345] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000001: edge_mask_reg_512p2[346] <= 1'b1;
 		default: edge_mask_reg_512p2[346] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010: edge_mask_reg_512p2[347] <= 1'b1;
 		default: edge_mask_reg_512p2[347] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110011,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110101,
11'b11001110110,
11'b11101010011,
11'b11101010100,
11'b11101010101,
11'b11101100011,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[348] <= 1'b1;
 		default: edge_mask_reg_512p2[348] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101000,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110011,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001000011,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110011,
11'b11001110101,
11'b11001110110: edge_mask_reg_512p2[349] <= 1'b1;
 		default: edge_mask_reg_512p2[349] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p2[350] <= 1'b1;
 		default: edge_mask_reg_512p2[350] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101001,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p2[351] <= 1'b1;
 		default: edge_mask_reg_512p2[351] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101010100,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p2[352] <= 1'b1;
 		default: edge_mask_reg_512p2[352] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p2[353] <= 1'b1;
 		default: edge_mask_reg_512p2[353] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010001000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[354] <= 1'b1;
 		default: edge_mask_reg_512p2[354] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000010,
11'b10010000011: edge_mask_reg_512p2[355] <= 1'b1;
 		default: edge_mask_reg_512p2[355] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010000,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111101000,
11'b1111101001,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101: edge_mask_reg_512p2[356] <= 1'b1;
 		default: edge_mask_reg_512p2[356] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[357] <= 1'b1;
 		default: edge_mask_reg_512p2[357] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110111000,
11'b1110111001,
11'b10010000010,
11'b10010000011,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101: edge_mask_reg_512p2[358] <= 1'b1;
 		default: edge_mask_reg_512p2[358] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b11010010010,
11'b11010010011,
11'b11010100010,
11'b11010100011: edge_mask_reg_512p2[359] <= 1'b1;
 		default: edge_mask_reg_512p2[359] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101100111,
11'b11101110100,
11'b11101110101,
11'b11101110110: edge_mask_reg_512p2[360] <= 1'b1;
 		default: edge_mask_reg_512p2[360] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000010,
11'b1010000011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1011101001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011: edge_mask_reg_512p2[361] <= 1'b1;
 		default: edge_mask_reg_512p2[361] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101100011,
11'b11101110010,
11'b11101110011,
11'b11101110100,
11'b11110000010,
11'b11110000011: edge_mask_reg_512p2[362] <= 1'b1;
 		default: edge_mask_reg_512p2[362] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111010000,
11'b10111010011: edge_mask_reg_512p2[363] <= 1'b1;
 		default: edge_mask_reg_512p2[363] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111010000,
11'b10111010011: edge_mask_reg_512p2[364] <= 1'b1;
 		default: edge_mask_reg_512p2[364] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111000001,
11'b10111010000,
11'b10111010001,
11'b10111010011: edge_mask_reg_512p2[365] <= 1'b1;
 		default: edge_mask_reg_512p2[365] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100: edge_mask_reg_512p2[366] <= 1'b1;
 		default: edge_mask_reg_512p2[366] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111000011,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111110011,
11'b10111110100: edge_mask_reg_512p2[367] <= 1'b1;
 		default: edge_mask_reg_512p2[367] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10011110110,
11'b10111000011,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110011,
11'b10111110100: edge_mask_reg_512p2[368] <= 1'b1;
 		default: edge_mask_reg_512p2[368] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10111000011,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110001,
11'b10111110010,
11'b10111110011,
11'b10111110100,
11'b10111110101: edge_mask_reg_512p2[369] <= 1'b1;
 		default: edge_mask_reg_512p2[369] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111000000,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111010000,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100011: edge_mask_reg_512p2[370] <= 1'b1;
 		default: edge_mask_reg_512p2[370] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000010,
11'b10011000011: edge_mask_reg_512p2[371] <= 1'b1;
 		default: edge_mask_reg_512p2[371] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100011000,
11'b1100011001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101: edge_mask_reg_512p2[372] <= 1'b1;
 		default: edge_mask_reg_512p2[372] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100011000,
11'b1100011001,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011001,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10101000001,
11'b10101000010,
11'b10101000011,
11'b10101000100: edge_mask_reg_512p2[373] <= 1'b1;
 		default: edge_mask_reg_512p2[373] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10010000000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[374] <= 1'b1;
 		default: edge_mask_reg_512p2[374] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10101100,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111001,
11'b1110111010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b10110110011,
11'b10110110100: edge_mask_reg_512p2[375] <= 1'b1;
 		default: edge_mask_reg_512p2[375] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011001,
11'b111011010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[376] <= 1'b1;
 		default: edge_mask_reg_512p2[376] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[377] <= 1'b1;
 		default: edge_mask_reg_512p2[377] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p2[378] <= 1'b1;
 		default: edge_mask_reg_512p2[378] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[379] <= 1'b1;
 		default: edge_mask_reg_512p2[379] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[380] <= 1'b1;
 		default: edge_mask_reg_512p2[380] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110011000,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[381] <= 1'b1;
 		default: edge_mask_reg_512p2[381] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[382] <= 1'b1;
 		default: edge_mask_reg_512p2[382] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[383] <= 1'b1;
 		default: edge_mask_reg_512p2[383] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[384] <= 1'b1;
 		default: edge_mask_reg_512p2[384] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[385] <= 1'b1;
 		default: edge_mask_reg_512p2[385] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001010000,
11'b10001010001: edge_mask_reg_512p2[386] <= 1'b1;
 		default: edge_mask_reg_512p2[386] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110101,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100011,
11'b10111100100,
11'b11011000001,
11'b11011000010: edge_mask_reg_512p2[387] <= 1'b1;
 		default: edge_mask_reg_512p2[387] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111000,
11'b1110111001,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010110101,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b11011000001,
11'b11011000010: edge_mask_reg_512p2[388] <= 1'b1;
 		default: edge_mask_reg_512p2[388] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111000,
11'b1110111001,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b10010110101,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110011,
11'b10111110100,
11'b11011000001,
11'b11011000010: edge_mask_reg_512p2[389] <= 1'b1;
 		default: edge_mask_reg_512p2[389] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11001011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b111011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111000,
11'b1110111001,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010110101,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b10111100010,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b11011000010,
11'b11011000011,
11'b11011010010,
11'b11011010011,
11'b11011010100,
11'b11011100010,
11'b11011100011,
11'b11011100100: edge_mask_reg_512p2[390] <= 1'b1;
 		default: edge_mask_reg_512p2[390] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100011,
11'b1111100100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100011,
11'b10011100100,
11'b10111000001,
11'b10111000010,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b11011000001,
11'b11011000010: edge_mask_reg_512p2[391] <= 1'b1;
 		default: edge_mask_reg_512p2[391] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100110,
11'b10110100111,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11110010011,
11'b11110010100: edge_mask_reg_512p2[392] <= 1'b1;
 		default: edge_mask_reg_512p2[392] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111011000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010010,
11'b10010010011,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[393] <= 1'b1;
 		default: edge_mask_reg_512p2[393] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1011011001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p2[394] <= 1'b1;
 		default: edge_mask_reg_512p2[394] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111001,
11'b101111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b11010100011,
11'b11010110011,
11'b11010110100: edge_mask_reg_512p2[395] <= 1'b1;
 		default: edge_mask_reg_512p2[395] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111001,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000011011,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b10000100110,
11'b10000100111,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000010,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b11000110010,
11'b11000110011,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000010,
11'b11001000011,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11100110100,
11'b11101000100: edge_mask_reg_512p2[396] <= 1'b1;
 		default: edge_mask_reg_512p2[396] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000010,
11'b10010000011: edge_mask_reg_512p2[397] <= 1'b1;
 		default: edge_mask_reg_512p2[397] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000001000,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101,
11'b11000000110,
11'b11000010011,
11'b11000010100,
11'b11000010101,
11'b11000010110,
11'b11100000010,
11'b11100000011,
11'b11100000100,
11'b11100000101,
11'b11100010011,
11'b11100010100,
11'b11100010101: edge_mask_reg_512p2[398] <= 1'b1;
 		default: edge_mask_reg_512p2[398] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010000001,
11'b10010010000: edge_mask_reg_512p2[399] <= 1'b1;
 		default: edge_mask_reg_512p2[399] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p2[400] <= 1'b1;
 		default: edge_mask_reg_512p2[400] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[401] <= 1'b1;
 		default: edge_mask_reg_512p2[401] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010010000: edge_mask_reg_512p2[402] <= 1'b1;
 		default: edge_mask_reg_512p2[402] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010000,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010000,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100111,
11'b1111101000: edge_mask_reg_512p2[403] <= 1'b1;
 		default: edge_mask_reg_512p2[403] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11001011,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110101010,
11'b10110111000,
11'b10110111001,
11'b10110111010,
11'b11010000111,
11'b11010001000,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010111000,
11'b11010111001,
11'b11110010101,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100101,
11'b11110100110,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p2[404] <= 1'b1;
 		default: edge_mask_reg_512p2[404] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100100100,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b10000110000,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100110001,
11'b10101000001,
11'b10101000010: edge_mask_reg_512p2[405] <= 1'b1;
 		default: edge_mask_reg_512p2[405] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b111011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100011000,
11'b1100011001,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101001,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100110001,
11'b10101000001,
11'b10101000010: edge_mask_reg_512p2[406] <= 1'b1;
 		default: edge_mask_reg_512p2[406] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101: edge_mask_reg_512p2[407] <= 1'b1;
 		default: edge_mask_reg_512p2[407] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100101,
11'b1100100110,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101: edge_mask_reg_512p2[408] <= 1'b1;
 		default: edge_mask_reg_512p2[408] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b11000000010,
11'b11000010010: edge_mask_reg_512p2[409] <= 1'b1;
 		default: edge_mask_reg_512p2[409] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111001,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b11000000010: edge_mask_reg_512p2[410] <= 1'b1;
 		default: edge_mask_reg_512p2[410] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b11000000001,
11'b11000000010,
11'b11000000011,
11'b11000000100: edge_mask_reg_512p2[411] <= 1'b1;
 		default: edge_mask_reg_512p2[411] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100010011,
11'b10100010100,
11'b11000000001,
11'b11000000010,
11'b11000000011,
11'b11000000100,
11'b11000000101: edge_mask_reg_512p2[412] <= 1'b1;
 		default: edge_mask_reg_512p2[412] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011001,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101010100,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p2[413] <= 1'b1;
 		default: edge_mask_reg_512p2[413] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p2[414] <= 1'b1;
 		default: edge_mask_reg_512p2[414] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110001,
11'b1110110010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b10010010000: edge_mask_reg_512p2[415] <= 1'b1;
 		default: edge_mask_reg_512p2[415] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110010,
11'b11101110011,
11'b11101110100,
11'b11110000010,
11'b11110000011: edge_mask_reg_512p2[416] <= 1'b1;
 		default: edge_mask_reg_512p2[416] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10011000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000110011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110010,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[417] <= 1'b1;
 		default: edge_mask_reg_512p2[417] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001: edge_mask_reg_512p2[418] <= 1'b1;
 		default: edge_mask_reg_512p2[418] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[419] <= 1'b1;
 		default: edge_mask_reg_512p2[419] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b1110101001,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011: edge_mask_reg_512p2[420] <= 1'b1;
 		default: edge_mask_reg_512p2[420] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101100011,
11'b1101100100,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b1110101001,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011: edge_mask_reg_512p2[421] <= 1'b1;
 		default: edge_mask_reg_512p2[421] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11110100011,
11'b11110100100,
11'b11110100101,
11'b11110110100,
11'b11110110101: edge_mask_reg_512p2[422] <= 1'b1;
 		default: edge_mask_reg_512p2[422] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b111011011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100011,
11'b1011100100,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111101000,
11'b1111101001,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100: edge_mask_reg_512p2[423] <= 1'b1;
 		default: edge_mask_reg_512p2[423] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[424] <= 1'b1;
 		default: edge_mask_reg_512p2[424] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000010,
11'b10010000011,
11'b10101100000,
11'b10101100001,
11'b10101100011: edge_mask_reg_512p2[425] <= 1'b1;
 		default: edge_mask_reg_512p2[425] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000010,
11'b10010000011,
11'b10101010000,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011: edge_mask_reg_512p2[426] <= 1'b1;
 		default: edge_mask_reg_512p2[426] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[427] <= 1'b1;
 		default: edge_mask_reg_512p2[427] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[428] <= 1'b1;
 		default: edge_mask_reg_512p2[428] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[429] <= 1'b1;
 		default: edge_mask_reg_512p2[429] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[430] <= 1'b1;
 		default: edge_mask_reg_512p2[430] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[431] <= 1'b1;
 		default: edge_mask_reg_512p2[431] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[432] <= 1'b1;
 		default: edge_mask_reg_512p2[432] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[433] <= 1'b1;
 		default: edge_mask_reg_512p2[433] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[434] <= 1'b1;
 		default: edge_mask_reg_512p2[434] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001100011,
11'b10001100100,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10101110001,
11'b10110000001: edge_mask_reg_512p2[435] <= 1'b1;
 		default: edge_mask_reg_512p2[435] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p2[436] <= 1'b1;
 		default: edge_mask_reg_512p2[436] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b10000000101,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100001,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110001,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100,
11'b10100010101,
11'b10100100001,
11'b10100100010,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110001,
11'b10100110010,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100: edge_mask_reg_512p2[437] <= 1'b1;
 		default: edge_mask_reg_512p2[437] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[438] <= 1'b1;
 		default: edge_mask_reg_512p2[438] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011000,
11'b1000011001: edge_mask_reg_512p2[439] <= 1'b1;
 		default: edge_mask_reg_512p2[439] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010011,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[440] <= 1'b1;
 		default: edge_mask_reg_512p2[440] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000111,
11'b1011001000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110110,
11'b1110110111,
11'b1110111000: edge_mask_reg_512p2[441] <= 1'b1;
 		default: edge_mask_reg_512p2[441] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110111,
11'b1010111000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010011,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[442] <= 1'b1;
 		default: edge_mask_reg_512p2[442] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010000,
11'b1000010001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000000,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010000,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000000000,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000010000,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10100000001,
11'b10100000010,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100: edge_mask_reg_512p2[443] <= 1'b1;
 		default: edge_mask_reg_512p2[443] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000001,
11'b110000010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000111,
11'b1111001000,
11'b10010010000,
11'b10010010010,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010110000,
11'b10010110001: edge_mask_reg_512p2[444] <= 1'b1;
 		default: edge_mask_reg_512p2[444] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101000,
11'b100101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1100011000,
11'b1100011001,
11'b10000000110,
11'b10100000100,
11'b10100000101,
11'b10100000110,
11'b10100000111,
11'b11000000100,
11'b11000000101,
11'b11000000110: edge_mask_reg_512p2[445] <= 1'b1;
 		default: edge_mask_reg_512p2[445] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10110000000,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100: edge_mask_reg_512p2[446] <= 1'b1;
 		default: edge_mask_reg_512p2[446] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000011,
11'b1000100,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b1101101000,
11'b1101101001,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p2[447] <= 1'b1;
 		default: edge_mask_reg_512p2[447] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[448] <= 1'b1;
 		default: edge_mask_reg_512p2[448] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110100000,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[449] <= 1'b1;
 		default: edge_mask_reg_512p2[449] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111011000,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110010,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p2[450] <= 1'b1;
 		default: edge_mask_reg_512p2[450] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10010000001: edge_mask_reg_512p2[451] <= 1'b1;
 		default: edge_mask_reg_512p2[451] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[452] <= 1'b1;
 		default: edge_mask_reg_512p2[452] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110010,
11'b10110011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101111000,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[453] <= 1'b1;
 		default: edge_mask_reg_512p2[453] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010010,
11'b1101010011,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[454] <= 1'b1;
 		default: edge_mask_reg_512p2[454] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[455] <= 1'b1;
 		default: edge_mask_reg_512p2[455] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110000,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010: edge_mask_reg_512p2[456] <= 1'b1;
 		default: edge_mask_reg_512p2[456] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100011,
11'b10101100100,
11'b10101110000,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p2[457] <= 1'b1;
 		default: edge_mask_reg_512p2[457] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p2[458] <= 1'b1;
 		default: edge_mask_reg_512p2[458] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100001000,
11'b1100001001,
11'b1100010001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000000111,
11'b10000010001,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010001,
11'b10100010010,
11'b10100010011,
11'b10100010100: edge_mask_reg_512p2[459] <= 1'b1;
 		default: edge_mask_reg_512p2[459] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[460] <= 1'b1;
 		default: edge_mask_reg_512p2[460] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110001000,
11'b110001001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010001000,
11'b1010001001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p2[461] <= 1'b1;
 		default: edge_mask_reg_512p2[461] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[462] <= 1'b1;
 		default: edge_mask_reg_512p2[462] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[463] <= 1'b1;
 		default: edge_mask_reg_512p2[463] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[464] <= 1'b1;
 		default: edge_mask_reg_512p2[464] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110000,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001: edge_mask_reg_512p2[465] <= 1'b1;
 		default: edge_mask_reg_512p2[465] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11000110,
11'b11000111,
11'b11001000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111110000,
11'b1111110001,
11'b1111110010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111100000,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111110000,
11'b10111110001,
11'b10111110010,
11'b10111110011: edge_mask_reg_512p2[466] <= 1'b1;
 		default: edge_mask_reg_512p2[466] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010110111,
11'b1010111000,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110000,
11'b1111110001,
11'b1111110010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011010000,
11'b10011010001,
11'b10011010010,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111010001,
11'b10111010010,
11'b10111010011,
11'b10111010100,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111110001,
11'b10111110010,
11'b10111110011: edge_mask_reg_512p2[467] <= 1'b1;
 		default: edge_mask_reg_512p2[467] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11000110,
11'b11000111,
11'b11001000,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1011000111,
11'b1011001000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100000,
11'b1111100001,
11'b1111100010,
11'b1111100011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110000,
11'b1111110001,
11'b1111110010,
11'b1111110011,
11'b1111110100,
11'b1111110101,
11'b1111110110,
11'b1111110111,
11'b1111111000,
11'b10011010011,
11'b10011100000,
11'b10011100001,
11'b10011100010,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011110000,
11'b10011110001,
11'b10011110010,
11'b10011110011,
11'b10011110100,
11'b10011110101,
11'b10111100001,
11'b10111100010,
11'b10111100011,
11'b10111110001,
11'b10111110010,
11'b10111110011: edge_mask_reg_512p2[468] <= 1'b1;
 		default: edge_mask_reg_512p2[468] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001: edge_mask_reg_512p2[469] <= 1'b1;
 		default: edge_mask_reg_512p2[469] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010010101,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110010,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000011,
11'b11011000100,
11'b11110100011,
11'b11110100100,
11'b11110100101,
11'b11110110011,
11'b11110110100,
11'b11110110101,
11'b11111000011,
11'b11111000100: edge_mask_reg_512p2[470] <= 1'b1;
 		default: edge_mask_reg_512p2[470] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p2[471] <= 1'b1;
 		default: edge_mask_reg_512p2[471] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110110,
11'b1110110111,
11'b1110111000: edge_mask_reg_512p2[472] <= 1'b1;
 		default: edge_mask_reg_512p2[472] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000: edge_mask_reg_512p2[473] <= 1'b1;
 		default: edge_mask_reg_512p2[473] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110111000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[474] <= 1'b1;
 		default: edge_mask_reg_512p2[474] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110111000,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p2[475] <= 1'b1;
 		default: edge_mask_reg_512p2[475] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001100010,
11'b11001100011,
11'b11001110010,
11'b11001110011: edge_mask_reg_512p2[476] <= 1'b1;
 		default: edge_mask_reg_512p2[476] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000010,
11'b10010000011,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[477] <= 1'b1;
 		default: edge_mask_reg_512p2[477] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010000,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010000,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100111,
11'b1111101000: edge_mask_reg_512p2[478] <= 1'b1;
 		default: edge_mask_reg_512p2[478] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001: edge_mask_reg_512p2[479] <= 1'b1;
 		default: edge_mask_reg_512p2[479] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b100100000,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010000,
11'b1000010001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100000,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100011000,
11'b1100011001,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101001000,
11'b1101001001: edge_mask_reg_512p2[480] <= 1'b1;
 		default: edge_mask_reg_512p2[480] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b100100000,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010000,
11'b1000010001,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000100000,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1100010010,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100000,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110000,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001: edge_mask_reg_512p2[481] <= 1'b1;
 		default: edge_mask_reg_512p2[481] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000: edge_mask_reg_512p2[482] <= 1'b1;
 		default: edge_mask_reg_512p2[482] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111011000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[483] <= 1'b1;
 		default: edge_mask_reg_512p2[483] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000111,
11'b1111001000,
11'b1111001001: edge_mask_reg_512p2[484] <= 1'b1;
 		default: edge_mask_reg_512p2[484] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001: edge_mask_reg_512p2[485] <= 1'b1;
 		default: edge_mask_reg_512p2[485] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000011010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100000001,
11'b1100000010,
11'b1100000011,
11'b1100000100,
11'b1100000101,
11'b1100000110,
11'b1100000111,
11'b1100010011,
11'b1100010100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101001,
11'b10000000001,
11'b10000000010,
11'b10000000011,
11'b10000000100,
11'b10000000101,
11'b10000000110,
11'b10000010010,
11'b10000010011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10100000001,
11'b10100000010,
11'b10100000011,
11'b10100000100,
11'b10100000101,
11'b10100010011,
11'b10100010100,
11'b10100010101: edge_mask_reg_512p2[486] <= 1'b1;
 		default: edge_mask_reg_512p2[486] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[487] <= 1'b1;
 		default: edge_mask_reg_512p2[487] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10011000000,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[488] <= 1'b1;
 		default: edge_mask_reg_512p2[488] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10110110001: edge_mask_reg_512p2[489] <= 1'b1;
 		default: edge_mask_reg_512p2[489] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10011000000,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[490] <= 1'b1;
 		default: edge_mask_reg_512p2[490] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010001000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010100010,
11'b10010100011,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10011000000,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p2[491] <= 1'b1;
 		default: edge_mask_reg_512p2[491] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110010,
11'b11110010011,
11'b11110010100,
11'b11110100010,
11'b11110100011,
11'b11110100100: edge_mask_reg_512p2[492] <= 1'b1;
 		default: edge_mask_reg_512p2[492] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100: edge_mask_reg_512p2[493] <= 1'b1;
 		default: edge_mask_reg_512p2[493] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100: edge_mask_reg_512p2[494] <= 1'b1;
 		default: edge_mask_reg_512p2[494] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p2[495] <= 1'b1;
 		default: edge_mask_reg_512p2[495] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11101010011,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101110011,
11'b11101110100,
11'b11101110101: edge_mask_reg_512p2[496] <= 1'b1;
 		default: edge_mask_reg_512p2[496] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100010,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p2[497] <= 1'b1;
 		default: edge_mask_reg_512p2[497] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110111000,
11'b1110111001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101: edge_mask_reg_512p2[498] <= 1'b1;
 		default: edge_mask_reg_512p2[498] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101000010,
11'b1101000011,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001: edge_mask_reg_512p2[499] <= 1'b1;
 		default: edge_mask_reg_512p2[499] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001: edge_mask_reg_512p2[500] <= 1'b1;
 		default: edge_mask_reg_512p2[500] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001: edge_mask_reg_512p2[501] <= 1'b1;
 		default: edge_mask_reg_512p2[501] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101000001,
11'b1101000010,
11'b1101000100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001: edge_mask_reg_512p2[502] <= 1'b1;
 		default: edge_mask_reg_512p2[502] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010000,
11'b10001010001,
11'b10001100000,
11'b10001100001: edge_mask_reg_512p2[503] <= 1'b1;
 		default: edge_mask_reg_512p2[503] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101011000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110010,
11'b10010000000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p2[504] <= 1'b1;
 		default: edge_mask_reg_512p2[504] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000000,
11'b10011000001,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101: edge_mask_reg_512p2[505] <= 1'b1;
 		default: edge_mask_reg_512p2[505] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010010,
11'b110010011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010000,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100010,
11'b1011100011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010000,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100111,
11'b1111101000,
11'b1111101001: edge_mask_reg_512p2[506] <= 1'b1;
 		default: edge_mask_reg_512p2[506] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010010,
11'b10010010011,
11'b10010100010,
11'b10010100011,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[507] <= 1'b1;
 		default: edge_mask_reg_512p2[507] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100010,
11'b10010100011,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[508] <= 1'b1;
 		default: edge_mask_reg_512p2[508] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010100010,
11'b10010100011,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p2[509] <= 1'b1;
 		default: edge_mask_reg_512p2[509] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p2[510] <= 1'b1;
 		default: edge_mask_reg_512p2[510] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p2[511] <= 1'b1;
 		default: edge_mask_reg_512p2[511] <= 1'b0;
 	endcase

end
endmodule

