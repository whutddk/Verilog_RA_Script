/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 7
date: 7
hour: 16
minutes: 35
second: 53
********************************************/

module prm_LUTX1chkp6(
	input [3:0] x,
	input [4:0] y,
	input [4:0] z,
	output [741:0] edge_mask_p6
);

	reg [741:0] edge_mask_reg_p6;
	assign edge_mask_p6= edge_mask_reg_p6;

always @( * ) begin
    case({z,y,x})
	14'b1010001100100,
	14'b1010001100101,
	14'b1010001100110,
	14'b1010001110100,
	14'b1010001110101,
	14'b1010001110110,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010000110,
	14'b1011001100100,
	14'b1011001100101,
	14'b1011001100110,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1100001100100,
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010101,
	14'b1101001010100,
	14'b1101001010101,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1110001010100,
	14'b1110001010101,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110011,
	14'b1110010110100,
	14'b1111001010100,
	14'b1111001010101,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001010100,
	14'b10000001010101,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[0] <= 1'b1;
 		default: edge_mask_reg_p6[0] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100101,
	14'b1010001100110,
	14'b1010001100111,
	14'b1010001110101,
	14'b1010001110110,
	14'b1010001110111,
	14'b1010010000101,
	14'b1010010000110,
	14'b1010010000111,
	14'b1011001100101,
	14'b1011001100110,
	14'b1011001100111,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010110,
	14'b1101001010101,
	14'b1101001010110,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1110001010101,
	14'b1110001010110,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001010101,
	14'b1111001010110,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000001010101,
	14'b10000001010110,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[1] <= 1'b1;
 		default: edge_mask_reg_p6[1] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100110,
	14'b1010001100111,
	14'b1010001101000,
	14'b1010001110110,
	14'b1010001110111,
	14'b1010001111000,
	14'b1010010000110,
	14'b1010010000111,
	14'b1010010001000,
	14'b1011001100110,
	14'b1011001100111,
	14'b1011001101000,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1101001010110,
	14'b1101001010111,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001010110,
	14'b1110001010111,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111001010110,
	14'b1111001010111,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010110,
	14'b10000001010111,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[2] <= 1'b1;
 		default: edge_mask_reg_p6[2] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100111,
	14'b1010001101000,
	14'b1010001101001,
	14'b1010001110111,
	14'b1010001111000,
	14'b1010001111001,
	14'b1010010000111,
	14'b1010010001000,
	14'b1010010001001,
	14'b1011001100111,
	14'b1011001101000,
	14'b1011001101001,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1101001010111,
	14'b1101001011000,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1110001010111,
	14'b1110001011000,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100000,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000001,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111001010111,
	14'b1111001011000,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b10000001010111,
	14'b10000001011000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[3] <= 1'b1;
 		default: edge_mask_reg_p6[3] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001101000,
	14'b1010001101001,
	14'b1010001101010,
	14'b1010001111000,
	14'b1010001111001,
	14'b1010001111010,
	14'b1010010001000,
	14'b1010010001001,
	14'b1010010001010,
	14'b1011001101000,
	14'b1011001101001,
	14'b1011001101010,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011001111010,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001101010,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101001011000,
	14'b1101001011001,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001101010,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101001111011,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010001011,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010011011,
	14'b1101010100000,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110001011000,
	14'b1110001011001,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001101010,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110001111011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010001011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1111001011000,
	14'b1111001011001,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001101010,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111001111011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001011000,
	14'b10000001011001,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001101010,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000001111011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010001: edge_mask_reg_p6[4] <= 1'b1;
 		default: edge_mask_reg_p6[4] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110000,
	14'b1001010000000,
	14'b1001010010000,
	14'b1010001110000,
	14'b1010010000000,
	14'b1010010010000,
	14'b1011001110000,
	14'b1011010000000,
	14'b1011010010000,
	14'b1100001110000,
	14'b1100010000000,
	14'b1100010010000,
	14'b1100010010001,
	14'b1101001110000,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010110000: edge_mask_reg_p6[5] <= 1'b1;
 		default: edge_mask_reg_p6[5] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110000,
	14'b1001001110001,
	14'b1001010000000,
	14'b1001010000001,
	14'b1001010010000,
	14'b1001010010001,
	14'b1010001110000,
	14'b1010001110001,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010010000,
	14'b1010010010001,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1101001100000,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1110001100000,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001011000000,
	14'b10010010110000: edge_mask_reg_p6[6] <= 1'b1;
 		default: edge_mask_reg_p6[6] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110000,
	14'b1001001110001,
	14'b1001001110010,
	14'b1001010000000,
	14'b1001010000001,
	14'b1001010000010,
	14'b1001010010000,
	14'b1001010010001,
	14'b1001010010010,
	14'b1010001110000,
	14'b1010001110001,
	14'b1010001110010,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100001,
	14'b1100010100010,
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110000,
	14'b1101010110001,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10100011110000: edge_mask_reg_p6[7] <= 1'b1;
 		default: edge_mask_reg_p6[7] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110001,
	14'b1001001110010,
	14'b1001001110011,
	14'b1001010000001,
	14'b1001010000010,
	14'b1001010000011,
	14'b1001010010001,
	14'b1001010010010,
	14'b1001010010011,
	14'b1010001110001,
	14'b1010001110010,
	14'b1010001110011,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100010,
	14'b1100010100011,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110001,
	14'b1101010110011,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10101011100000: edge_mask_reg_p6[8] <= 1'b1;
 		default: edge_mask_reg_p6[8] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110010,
	14'b1001001110011,
	14'b1001001110100,
	14'b1001010000010,
	14'b1001010000011,
	14'b1001010000100,
	14'b1001010010010,
	14'b1001010010011,
	14'b1001010010100,
	14'b1010001110010,
	14'b1010001110011,
	14'b1010001110100,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011001110100,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100011,
	14'b1100010100100,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[9] <= 1'b1;
 		default: edge_mask_reg_p6[9] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110011,
	14'b1001001110100,
	14'b1001001110101,
	14'b1001010000011,
	14'b1001010000100,
	14'b1001010000101,
	14'b1001010010011,
	14'b1001010010100,
	14'b1001010010101,
	14'b1010001110011,
	14'b1010001110100,
	14'b1010001110101,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010010101,
	14'b1011001110011,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100100,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[10] <= 1'b1;
 		default: edge_mask_reg_p6[10] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001001110100,
	14'b1001001110101,
	14'b1001001110110,
	14'b1001010000100,
	14'b1001010000101,
	14'b1001010000110,
	14'b1001010010100,
	14'b1001010010101,
	14'b1001010010110,
	14'b1010001110100,
	14'b1010001110101,
	14'b1010001110110,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010000110,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010010110,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100101,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[11] <= 1'b1;
 		default: edge_mask_reg_p6[11] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110101,
	14'b1010001110110,
	14'b1010001110111,
	14'b1010010000101,
	14'b1010010000110,
	14'b1010010000111,
	14'b1010010010101,
	14'b1010010010110,
	14'b1010010010111,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100110,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000100,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010010000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[12] <= 1'b1;
 		default: edge_mask_reg_p6[12] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110110,
	14'b1010001110111,
	14'b1010001111000,
	14'b1010010000110,
	14'b1010010000111,
	14'b1010010001000,
	14'b1010010010110,
	14'b1010010010111,
	14'b1010010011000,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100111,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010000,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[13] <= 1'b1;
 		default: edge_mask_reg_p6[13] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110111,
	14'b1010001111000,
	14'b1010001111001,
	14'b1010010000111,
	14'b1010010001000,
	14'b1010010001001,
	14'b1010010010111,
	14'b1010010011000,
	14'b1010010011001,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010101000,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010: edge_mask_reg_p6[14] <= 1'b1;
 		default: edge_mask_reg_p6[14] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001111000,
	14'b1010001111001,
	14'b1010001111010,
	14'b1010010001000,
	14'b1010010001001,
	14'b1010010001010,
	14'b1010010011000,
	14'b1010010011001,
	14'b1010010011010,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011001111010,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101001,
	14'b1100011100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010001011,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010011011,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010101011,
	14'b1101010110000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010001011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010: edge_mask_reg_p6[15] <= 1'b1;
 		default: edge_mask_reg_p6[15] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000000,
	14'b1001010010000,
	14'b1001010100000,
	14'b1010010000000,
	14'b1010010010000,
	14'b1010010100000,
	14'b1011010000000,
	14'b1011010010000,
	14'b1011010100000,
	14'b1100010000000,
	14'b1100010010000,
	14'b1100010100000,
	14'b1100010100001,
	14'b1101010000000,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001010100000,
	14'b10001010110000: edge_mask_reg_p6[16] <= 1'b1;
 		default: edge_mask_reg_p6[16] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000000,
	14'b1001010000001,
	14'b1001010010000,
	14'b1001010010001,
	14'b1001010100000,
	14'b1001010100001,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010100000,
	14'b1010010100001,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1101001110000,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010011000000: edge_mask_reg_p6[17] <= 1'b1;
 		default: edge_mask_reg_p6[17] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000000,
	14'b1001010000001,
	14'b1001010000010,
	14'b1001010010000,
	14'b1001010010001,
	14'b1001010010010,
	14'b1001010100000,
	14'b1001010100001,
	14'b1001010100010,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110001,
	14'b1100010110010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011010000: edge_mask_reg_p6[18] <= 1'b1;
 		default: edge_mask_reg_p6[18] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000001,
	14'b1001010000010,
	14'b1001010000011,
	14'b1001010010001,
	14'b1001010010010,
	14'b1001010010011,
	14'b1001010100001,
	14'b1001010100010,
	14'b1001010100011,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110010,
	14'b1100010110011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[19] <= 1'b1;
 		default: edge_mask_reg_p6[19] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000010,
	14'b1001010000011,
	14'b1001010000100,
	14'b1001010010010,
	14'b1001010010011,
	14'b1001010010100,
	14'b1001010100010,
	14'b1001010100011,
	14'b1001010100100,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110011,
	14'b1100010110100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[20] <= 1'b1;
 		default: edge_mask_reg_p6[20] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000011,
	14'b1001010000100,
	14'b1001010000101,
	14'b1001010010011,
	14'b1001010010100,
	14'b1001010010101,
	14'b1001010100011,
	14'b1001010100100,
	14'b1001010100101,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110100,
	14'b1100010110101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011110000,
	14'b10001010000010,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[21] <= 1'b1;
 		default: edge_mask_reg_p6[21] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000100,
	14'b1001010000101,
	14'b1001010000110,
	14'b1001010010100,
	14'b1001010010101,
	14'b1001010010110,
	14'b1001010100100,
	14'b1001010100101,
	14'b1001010100110,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010000110,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010010110,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010100110,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110101,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000100,
	14'b1101011000101,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011110000,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010000011,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[22] <= 1'b1;
 		default: edge_mask_reg_p6[22] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010000101,
	14'b1001010000110,
	14'b1001010000111,
	14'b1001010010101,
	14'b1001010010110,
	14'b1001010010111,
	14'b1001010100101,
	14'b1001010100110,
	14'b1001010100111,
	14'b1010010000101,
	14'b1010010000110,
	14'b1010010000111,
	14'b1010010010101,
	14'b1010010010110,
	14'b1010010010111,
	14'b1010010100101,
	14'b1010010100110,
	14'b1010010100111,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110110,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10001010000100,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[23] <= 1'b1;
 		default: edge_mask_reg_p6[23] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000110,
	14'b1010010000111,
	14'b1010010001000,
	14'b1010010010110,
	14'b1010010010111,
	14'b1010010011000,
	14'b1010010100110,
	14'b1010010100111,
	14'b1010010101000,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110111,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010000101,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[24] <= 1'b1;
 		default: edge_mask_reg_p6[24] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000111,
	14'b1010010001000,
	14'b1010010001001,
	14'b1010010010111,
	14'b1010010011000,
	14'b1010010011001,
	14'b1010010100111,
	14'b1010010101000,
	14'b1010010101001,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010111000,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[25] <= 1'b1;
 		default: edge_mask_reg_p6[25] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010001000,
	14'b1010010001001,
	14'b1010010001010,
	14'b1010010011000,
	14'b1010010011001,
	14'b1010010011010,
	14'b1010010101000,
	14'b1010010101001,
	14'b1010010101010,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111001,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010011011,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010101011,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101010111011,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100001: edge_mask_reg_p6[26] <= 1'b1;
 		default: edge_mask_reg_p6[26] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010000,
	14'b1001010100000,
	14'b1001010110000,
	14'b1010010010000,
	14'b1010010100000,
	14'b1010010110000,
	14'b1011010010000,
	14'b1011010100000,
	14'b1011010110000,
	14'b1100010010000,
	14'b1100010100000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10001011000000: edge_mask_reg_p6[27] <= 1'b1;
 		default: edge_mask_reg_p6[27] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010000,
	14'b1001010010001,
	14'b1001010100000,
	14'b1001010100001,
	14'b1001010110000,
	14'b1001010110001,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010110000,
	14'b1010010110001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1101010000000,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010001,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011010000: edge_mask_reg_p6[28] <= 1'b1;
 		default: edge_mask_reg_p6[28] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010000,
	14'b1001010010001,
	14'b1001010010010,
	14'b1001010100000,
	14'b1001010100001,
	14'b1001010100010,
	14'b1001010110000,
	14'b1001010110001,
	14'b1001010110010,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000001,
	14'b1100011000010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10010011000000,
	14'b10010011010000: edge_mask_reg_p6[29] <= 1'b1;
 		default: edge_mask_reg_p6[29] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010001,
	14'b1001010010010,
	14'b1001010010011,
	14'b1001010100001,
	14'b1001010100010,
	14'b1001010100011,
	14'b1001010110001,
	14'b1001010110010,
	14'b1001010110011,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000010,
	14'b1100011000011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000: edge_mask_reg_p6[30] <= 1'b1;
 		default: edge_mask_reg_p6[30] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010010,
	14'b1001010010011,
	14'b1001010010100,
	14'b1001010100010,
	14'b1001010100011,
	14'b1001010100100,
	14'b1001010110010,
	14'b1001010110011,
	14'b1001010110100,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000011,
	14'b1100011000100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[31] <= 1'b1;
 		default: edge_mask_reg_p6[31] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010011,
	14'b1001010010100,
	14'b1001010010101,
	14'b1001010100011,
	14'b1001010100100,
	14'b1001010100101,
	14'b1001010110011,
	14'b1001010110100,
	14'b1001010110101,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000100,
	14'b1100011000101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100001,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[32] <= 1'b1;
 		default: edge_mask_reg_p6[32] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010100,
	14'b1001010010101,
	14'b1001010010110,
	14'b1001010100100,
	14'b1001010100101,
	14'b1001010100110,
	14'b1001010110100,
	14'b1001010110101,
	14'b1001010110110,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010010110,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010100110,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010010110110,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000101,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[33] <= 1'b1;
 		default: edge_mask_reg_p6[33] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010010101,
	14'b1001010010110,
	14'b1001010010111,
	14'b1001010100101,
	14'b1001010100110,
	14'b1001010100111,
	14'b1001010110101,
	14'b1001010110110,
	14'b1001010110111,
	14'b1010010010101,
	14'b1010010010110,
	14'b1010010010111,
	14'b1010010100101,
	14'b1010010100110,
	14'b1010010100111,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010010110111,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000110,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010101,
	14'b1101011010110,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010100000,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[34] <= 1'b1;
 		default: edge_mask_reg_p6[34] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010110,
	14'b1010010010111,
	14'b1010010011000,
	14'b1010010100110,
	14'b1010010100111,
	14'b1010010101000,
	14'b1010010110110,
	14'b1010010110111,
	14'b1010010111000,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000111,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010110,
	14'b1101011010111,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[35] <= 1'b1;
 		default: edge_mask_reg_p6[35] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010111,
	14'b1010010011000,
	14'b1010010011001,
	14'b1010010100111,
	14'b1010010101000,
	14'b1010010101001,
	14'b1010010110111,
	14'b1010010111000,
	14'b1010010111001,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011001000,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101100000000,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[36] <= 1'b1;
 		default: edge_mask_reg_p6[36] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010011000,
	14'b1010010011001,
	14'b1010010011010,
	14'b1010010101000,
	14'b1010010101001,
	14'b1010010101010,
	14'b1010010111000,
	14'b1010010111001,
	14'b1010010111010,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001001,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010101011,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101010111011,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011001011,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010: edge_mask_reg_p6[37] <= 1'b1;
 		default: edge_mask_reg_p6[37] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100000,
	14'b1001010110000,
	14'b1001011000000,
	14'b1010010100000,
	14'b1010010110000,
	14'b1010011000000,
	14'b1011010100000,
	14'b1011010110000,
	14'b1011011000000,
	14'b1100010100000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001: edge_mask_reg_p6[38] <= 1'b1;
 		default: edge_mask_reg_p6[38] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100000,
	14'b1001010100001,
	14'b1001010110000,
	14'b1001010110001,
	14'b1001011000000,
	14'b1001011000001,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010011000000,
	14'b1010011000001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1101010010000,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10001011010000,
	14'b10001011100000: edge_mask_reg_p6[39] <= 1'b1;
 		default: edge_mask_reg_p6[39] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100000,
	14'b1001010100001,
	14'b1001010100010,
	14'b1001010110000,
	14'b1001010110001,
	14'b1001010110010,
	14'b1001011000000,
	14'b1001011000001,
	14'b1001011000010,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010001,
	14'b1100011010010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010011010000,
	14'b10010011100000: edge_mask_reg_p6[40] <= 1'b1;
 		default: edge_mask_reg_p6[40] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100001,
	14'b1001010100010,
	14'b1001010100011,
	14'b1001010110001,
	14'b1001010110010,
	14'b1001010110011,
	14'b1001011000001,
	14'b1001011000010,
	14'b1001011000011,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001: edge_mask_reg_p6[41] <= 1'b1;
 		default: edge_mask_reg_p6[41] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100010,
	14'b1001010100011,
	14'b1001010100100,
	14'b1001010110010,
	14'b1001010110011,
	14'b1001010110100,
	14'b1001011000010,
	14'b1001011000011,
	14'b1001011000100,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100100000000: edge_mask_reg_p6[42] <= 1'b1;
 		default: edge_mask_reg_p6[42] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100011,
	14'b1001010100100,
	14'b1001010100101,
	14'b1001010110011,
	14'b1001010110100,
	14'b1001010110101,
	14'b1001011000011,
	14'b1001011000100,
	14'b1001011000101,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[43] <= 1'b1;
 		default: edge_mask_reg_p6[43] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100100,
	14'b1001010100101,
	14'b1001010100110,
	14'b1001010110100,
	14'b1001010110101,
	14'b1001010110110,
	14'b1001011000100,
	14'b1001011000101,
	14'b1001011000110,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010100110,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011000110,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000100000000,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[44] <= 1'b1;
 		default: edge_mask_reg_p6[44] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100101,
	14'b1001010100110,
	14'b1001010100111,
	14'b1001010110101,
	14'b1001010110110,
	14'b1001010110111,
	14'b1001011000101,
	14'b1001011000110,
	14'b1001011000111,
	14'b1010010100101,
	14'b1010010100110,
	14'b1010010100111,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010010110111,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011000111,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111100000000,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010110000,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000: edge_mask_reg_p6[45] <= 1'b1;
 		default: edge_mask_reg_p6[45] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010100110,
	14'b1001010100111,
	14'b1001010101000,
	14'b1001010110110,
	14'b1001010110111,
	14'b1001010111000,
	14'b1001011000110,
	14'b1001011000111,
	14'b1001011001000,
	14'b1010010100110,
	14'b1010010100111,
	14'b1010010101000,
	14'b1010010110110,
	14'b1010010110111,
	14'b1010010111000,
	14'b1010011000110,
	14'b1010011000111,
	14'b1010011001000,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000: edge_mask_reg_p6[46] <= 1'b1;
 		default: edge_mask_reg_p6[46] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100111,
	14'b1010010101000,
	14'b1010010101001,
	14'b1010010110111,
	14'b1010010111000,
	14'b1010010111001,
	14'b1010011000111,
	14'b1010011001000,
	14'b1010011001001,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011011000,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011100111,
	14'b1101011101000,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000: edge_mask_reg_p6[47] <= 1'b1;
 		default: edge_mask_reg_p6[47] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010101000,
	14'b1010010101001,
	14'b1010010101010,
	14'b1010010111000,
	14'b1010010111001,
	14'b1010010111010,
	14'b1010011001000,
	14'b1010011001001,
	14'b1010011001010,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011001,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101010111011,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011001011,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011011011,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100001,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110001: edge_mask_reg_p6[48] <= 1'b1;
 		default: edge_mask_reg_p6[48] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110000,
	14'b1001011000000,
	14'b1001011010000,
	14'b1010010110000,
	14'b1010011000000,
	14'b1010011010000,
	14'b1011010110000,
	14'b1011011000000,
	14'b1011011010000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001: edge_mask_reg_p6[49] <= 1'b1;
 		default: edge_mask_reg_p6[49] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110000,
	14'b1001010110001,
	14'b1001011000000,
	14'b1001011000001,
	14'b1001011010000,
	14'b1001011010001,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011010000,
	14'b1010011010001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001011100000,
	14'b10001011110000: edge_mask_reg_p6[50] <= 1'b1;
 		default: edge_mask_reg_p6[50] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110000,
	14'b1001010110001,
	14'b1001010110010,
	14'b1001011000000,
	14'b1001011000001,
	14'b1001011000010,
	14'b1001011010000,
	14'b1001011010001,
	14'b1001011010010,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010011100000,
	14'b10010011110000: edge_mask_reg_p6[51] <= 1'b1;
 		default: edge_mask_reg_p6[51] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110001,
	14'b1001010110010,
	14'b1001010110011,
	14'b1001011000001,
	14'b1001011000010,
	14'b1001011000011,
	14'b1001011010001,
	14'b1001011010010,
	14'b1001011010011,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001: edge_mask_reg_p6[52] <= 1'b1;
 		default: edge_mask_reg_p6[52] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110010,
	14'b1001010110011,
	14'b1001010110100,
	14'b1001011000010,
	14'b1001011000011,
	14'b1001011000100,
	14'b1001011010010,
	14'b1001011010011,
	14'b1001011010100,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000: edge_mask_reg_p6[53] <= 1'b1;
 		default: edge_mask_reg_p6[53] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110011,
	14'b1001010110100,
	14'b1001010110101,
	14'b1001011000011,
	14'b1001011000100,
	14'b1001011000101,
	14'b1001011010011,
	14'b1001011010100,
	14'b1001011010101,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110011,
	14'b1101011110100,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[54] <= 1'b1;
 		default: edge_mask_reg_p6[54] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110100,
	14'b1001010110101,
	14'b1001010110110,
	14'b1001011000100,
	14'b1001011000101,
	14'b1001011000110,
	14'b1001011010100,
	14'b1001011010101,
	14'b1001011010110,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110100,
	14'b1101011110101,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[55] <= 1'b1;
 		default: edge_mask_reg_p6[55] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110101,
	14'b1001010110110,
	14'b1001010110111,
	14'b1001011000101,
	14'b1001011000110,
	14'b1001011000111,
	14'b1001011010101,
	14'b1001011010110,
	14'b1001011010111,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010010110111,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011000111,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011010111,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110101,
	14'b1101011110110,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[56] <= 1'b1;
 		default: edge_mask_reg_p6[56] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001010110110,
	14'b1001010110111,
	14'b1001010111000,
	14'b1001011000110,
	14'b1001011000111,
	14'b1001011001000,
	14'b1001011010110,
	14'b1001011010111,
	14'b1001011011000,
	14'b1010010110110,
	14'b1010010110111,
	14'b1010010111000,
	14'b1010011000110,
	14'b1010011000111,
	14'b1010011001000,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011011000,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110110,
	14'b1101011110111,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[57] <= 1'b1;
 		default: edge_mask_reg_p6[57] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110111,
	14'b1010010111000,
	14'b1010010111001,
	14'b1010011000111,
	14'b1010011001000,
	14'b1010011001001,
	14'b1010011010111,
	14'b1010011011000,
	14'b1010011011001,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011110111,
	14'b1101011111000,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[58] <= 1'b1;
 		default: edge_mask_reg_p6[58] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010111000,
	14'b1010010111001,
	14'b1010010111010,
	14'b1010011001000,
	14'b1010011001001,
	14'b1010011001010,
	14'b1010011011000,
	14'b1010011011001,
	14'b1010011011010,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101001,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011001011,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011011011,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011101011,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000000,
	14'b1101100010000,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010000,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010: edge_mask_reg_p6[59] <= 1'b1;
 		default: edge_mask_reg_p6[59] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000000,
	14'b1001011010000,
	14'b1001011100000,
	14'b1010011000000,
	14'b1010011010000,
	14'b1010011100000,
	14'b1011011000000,
	14'b1011011010000,
	14'b1011011100000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001: edge_mask_reg_p6[60] <= 1'b1;
 		default: edge_mask_reg_p6[60] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000000,
	14'b1001011000001,
	14'b1001011010000,
	14'b1001011010001,
	14'b1001011100000,
	14'b1001011100001,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011100000,
	14'b1010011100001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1101010110000,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10001011110000: edge_mask_reg_p6[61] <= 1'b1;
 		default: edge_mask_reg_p6[61] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000000,
	14'b1001011000001,
	14'b1001011000010,
	14'b1001011010000,
	14'b1001011010001,
	14'b1001011010010,
	14'b1001011100000,
	14'b1001011100001,
	14'b1001011100010,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000: edge_mask_reg_p6[62] <= 1'b1;
 		default: edge_mask_reg_p6[62] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000001,
	14'b1001011000010,
	14'b1001011000011,
	14'b1001011010001,
	14'b1001011010010,
	14'b1001011010011,
	14'b1001011100001,
	14'b1001011100010,
	14'b1001011100011,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000001,
	14'b1101100000010,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000: edge_mask_reg_p6[63] <= 1'b1;
 		default: edge_mask_reg_p6[63] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000010,
	14'b1001011000011,
	14'b1001011000100,
	14'b1001011010010,
	14'b1001011010011,
	14'b1001011010100,
	14'b1001011100010,
	14'b1001011100011,
	14'b1001011100100,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000010,
	14'b1101100000011,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011011100000,
	14'b10011011110000: edge_mask_reg_p6[64] <= 1'b1;
 		default: edge_mask_reg_p6[64] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000011,
	14'b1001011000100,
	14'b1001011000101,
	14'b1001011010011,
	14'b1001011010100,
	14'b1001011010101,
	14'b1001011100011,
	14'b1001011100100,
	14'b1001011100101,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000011,
	14'b1101100000100,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[65] <= 1'b1;
 		default: edge_mask_reg_p6[65] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000100,
	14'b1001011000101,
	14'b1001011000110,
	14'b1001011010100,
	14'b1001011010101,
	14'b1001011010110,
	14'b1001011100100,
	14'b1001011100101,
	14'b1001011100110,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[66] <= 1'b1;
 		default: edge_mask_reg_p6[66] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000101,
	14'b1001011000110,
	14'b1001011000111,
	14'b1001011010101,
	14'b1001011010110,
	14'b1001011010111,
	14'b1001011100101,
	14'b1001011100110,
	14'b1001011100111,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011000111,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011100111,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10001011000000,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10010011000000,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[67] <= 1'b1;
 		default: edge_mask_reg_p6[67] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011000110,
	14'b1001011000111,
	14'b1001011001000,
	14'b1001011010110,
	14'b1001011010111,
	14'b1001011011000,
	14'b1001011100110,
	14'b1001011100111,
	14'b1001011101000,
	14'b1010011000110,
	14'b1010011000111,
	14'b1010011001000,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011011000,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011101000,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010000,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[68] <= 1'b1;
 		default: edge_mask_reg_p6[68] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000111,
	14'b1010011001000,
	14'b1010011001001,
	14'b1010011010111,
	14'b1010011011000,
	14'b1010011011001,
	14'b1010011100111,
	14'b1010011101000,
	14'b1010011101001,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000000,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010000,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000: edge_mask_reg_p6[69] <= 1'b1;
 		default: edge_mask_reg_p6[69] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011001000,
	14'b1010011001001,
	14'b1010011001010,
	14'b1010011011000,
	14'b1010011011001,
	14'b1010011011010,
	14'b1010011101000,
	14'b1010011101001,
	14'b1010011101010,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011011011,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011101011,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100010000,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000000,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010000,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001: edge_mask_reg_p6[70] <= 1'b1;
 		default: edge_mask_reg_p6[70] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010000,
	14'b1001011100000,
	14'b1001011110000,
	14'b1010011010000,
	14'b1010011100000,
	14'b1010011110000,
	14'b1011011010000,
	14'b1011011100000,
	14'b1011011110000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000: edge_mask_reg_p6[71] <= 1'b1;
 		default: edge_mask_reg_p6[71] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010000,
	14'b1001011010001,
	14'b1001011100000,
	14'b1001011100001,
	14'b1001011110000,
	14'b1001011110001,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011110000,
	14'b1010011110001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001100000000: edge_mask_reg_p6[72] <= 1'b1;
 		default: edge_mask_reg_p6[72] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010000,
	14'b1001011010001,
	14'b1001011010010,
	14'b1001011100000,
	14'b1001011100001,
	14'b1001011100010,
	14'b1001011110000,
	14'b1001011110001,
	14'b1001011110010,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001: edge_mask_reg_p6[73] <= 1'b1;
 		default: edge_mask_reg_p6[73] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010001,
	14'b1001011010010,
	14'b1001011010011,
	14'b1001011100001,
	14'b1001011100010,
	14'b1001011100011,
	14'b1001011110001,
	14'b1001011110010,
	14'b1001011110011,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000: edge_mask_reg_p6[74] <= 1'b1;
 		default: edge_mask_reg_p6[74] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010010,
	14'b1001011010011,
	14'b1001011010100,
	14'b1001011100010,
	14'b1001011100011,
	14'b1001011100100,
	14'b1001011110010,
	14'b1001011110011,
	14'b1001011110100,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011011100000,
	14'b10011011110000: edge_mask_reg_p6[75] <= 1'b1;
 		default: edge_mask_reg_p6[75] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010011,
	14'b1001011010100,
	14'b1001011010101,
	14'b1001011100011,
	14'b1001011100100,
	14'b1001011100101,
	14'b1001011110011,
	14'b1001011110100,
	14'b1001011110101,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[76] <= 1'b1;
 		default: edge_mask_reg_p6[76] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010100,
	14'b1001011010101,
	14'b1001011010110,
	14'b1001011100100,
	14'b1001011100101,
	14'b1001011100110,
	14'b1001011110100,
	14'b1001011110101,
	14'b1001011110110,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[77] <= 1'b1;
 		default: edge_mask_reg_p6[77] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010101,
	14'b1001011010110,
	14'b1001011010111,
	14'b1001011100101,
	14'b1001011100110,
	14'b1001011100111,
	14'b1001011110101,
	14'b1001011110110,
	14'b1001011110111,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[78] <= 1'b1;
 		default: edge_mask_reg_p6[78] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011010110,
	14'b1001011010111,
	14'b1001011011000,
	14'b1001011100110,
	14'b1001011100111,
	14'b1001011101000,
	14'b1001011110110,
	14'b1001011110111,
	14'b1001011111000,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011011000,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011101000,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010011111000,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b10000011000000,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[79] <= 1'b1;
 		default: edge_mask_reg_p6[79] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010111,
	14'b1010011011000,
	14'b1010011011001,
	14'b1010011100111,
	14'b1010011101000,
	14'b1010011101001,
	14'b1010011110111,
	14'b1010011111000,
	14'b1010011111001,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1111011000000,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100000010: edge_mask_reg_p6[80] <= 1'b1;
 		default: edge_mask_reg_p6[80] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011011000,
	14'b1010011011001,
	14'b1010011011010,
	14'b1010011101000,
	14'b1010011101001,
	14'b1010011101010,
	14'b1010011111000,
	14'b1010011111001,
	14'b1010011111010,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011101011,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101011111011,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1110011000000,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010000,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100000,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000000,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011110001,
	14'b10101100000001: edge_mask_reg_p6[81] <= 1'b1;
 		default: edge_mask_reg_p6[81] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100000,
	14'b1001011110000,
	14'b1001100000000,
	14'b1010011100000,
	14'b1010011110000,
	14'b1010100000000,
	14'b1011011100000,
	14'b1011011110000,
	14'b1011100000000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100100000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100100000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000: edge_mask_reg_p6[82] <= 1'b1;
 		default: edge_mask_reg_p6[82] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100000,
	14'b1001011100001,
	14'b1001011110000,
	14'b1001011110001,
	14'b1001100000000,
	14'b1001100000001,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010100000000,
	14'b1010100000001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011100000000,
	14'b1011100000001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001: edge_mask_reg_p6[83] <= 1'b1;
 		default: edge_mask_reg_p6[83] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100000,
	14'b1001011100001,
	14'b1001011100010,
	14'b1001011110000,
	14'b1001011110001,
	14'b1001011110010,
	14'b1001100000000,
	14'b1001100000001,
	14'b1001100000010,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100000010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100000010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000: edge_mask_reg_p6[84] <= 1'b1;
 		default: edge_mask_reg_p6[84] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100001,
	14'b1001011100010,
	14'b1001011100011,
	14'b1001011110001,
	14'b1001011110010,
	14'b1001011110011,
	14'b1001100000001,
	14'b1001100000010,
	14'b1001100000011,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100000011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100000011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000: edge_mask_reg_p6[85] <= 1'b1;
 		default: edge_mask_reg_p6[85] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100010,
	14'b1001011100011,
	14'b1001011100100,
	14'b1001011110010,
	14'b1001011110011,
	14'b1001011110100,
	14'b1001100000010,
	14'b1001100000011,
	14'b1001100000100,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[86] <= 1'b1;
 		default: edge_mask_reg_p6[86] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100011,
	14'b1001011100100,
	14'b1001011100101,
	14'b1001011110011,
	14'b1001011110100,
	14'b1001011110101,
	14'b1001100000011,
	14'b1001100000100,
	14'b1001100000101,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000: edge_mask_reg_p6[87] <= 1'b1;
 		default: edge_mask_reg_p6[87] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100100,
	14'b1001011100101,
	14'b1001011100110,
	14'b1001011110100,
	14'b1001011110101,
	14'b1001011110110,
	14'b1001100000100,
	14'b1001100000101,
	14'b1001100000110,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[88] <= 1'b1;
 		default: edge_mask_reg_p6[88] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100101,
	14'b1001011100110,
	14'b1001011100111,
	14'b1001011110101,
	14'b1001011110110,
	14'b1001011110111,
	14'b1001100000101,
	14'b1001100000110,
	14'b1001100000111,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100000111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[89] <= 1'b1;
 		default: edge_mask_reg_p6[89] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011100110,
	14'b1001011100111,
	14'b1001011101000,
	14'b1001011110110,
	14'b1001011110111,
	14'b1001011111000,
	14'b1001100000110,
	14'b1001100000111,
	14'b1001100001000,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011101000,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010011111000,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100001000,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b10000011010000,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[90] <= 1'b1;
 		default: edge_mask_reg_p6[90] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100111,
	14'b1010011101000,
	14'b1010011101001,
	14'b1010011110111,
	14'b1010011111000,
	14'b1010011111001,
	14'b1010100000111,
	14'b1010100001000,
	14'b1010100001001,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1111011010000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100000,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101011110010,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100000010: edge_mask_reg_p6[91] <= 1'b1;
 		default: edge_mask_reg_p6[91] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011101000,
	14'b1010011101001,
	14'b1010011101010,
	14'b1010011111000,
	14'b1010011111001,
	14'b1010011111010,
	14'b1010100001000,
	14'b1010100001001,
	14'b1010100001010,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011101011,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101011111011,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100001011,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1110011010000,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100001011,
	14'b1110100010000,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[92] <= 1'b1;
 		default: edge_mask_reg_p6[92] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110000,
	14'b1001100000000,
	14'b1001100010000,
	14'b1010011110000,
	14'b1010100000000,
	14'b1010100010000,
	14'b1010100100000,
	14'b1011011110000,
	14'b1011100000000,
	14'b1011100010000,
	14'b1011100100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100110000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100110000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100110000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000: edge_mask_reg_p6[93] <= 1'b1;
 		default: edge_mask_reg_p6[93] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110000,
	14'b1001011110001,
	14'b1001100000000,
	14'b1001100000001,
	14'b1001100010000,
	14'b1001100010001,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100010000,
	14'b1010100010001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100010000,
	14'b1011100010001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10001011110000: edge_mask_reg_p6[94] <= 1'b1;
 		default: edge_mask_reg_p6[94] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110000,
	14'b1001011110001,
	14'b1001011110010,
	14'b1001100000000,
	14'b1001100000001,
	14'b1001100000010,
	14'b1001100010000,
	14'b1001100010001,
	14'b1001100010010,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100010010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100010010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000: edge_mask_reg_p6[95] <= 1'b1;
 		default: edge_mask_reg_p6[95] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110001,
	14'b1001011110010,
	14'b1001011110011,
	14'b1001100000001,
	14'b1001100000010,
	14'b1001100000011,
	14'b1001100010001,
	14'b1001100010010,
	14'b1001100010011,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100010011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100010011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[96] <= 1'b1;
 		default: edge_mask_reg_p6[96] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110010,
	14'b1001011110011,
	14'b1001011110100,
	14'b1001100000010,
	14'b1001100000011,
	14'b1001100000100,
	14'b1001100010010,
	14'b1001100010011,
	14'b1001100010100,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100010100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100010100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[97] <= 1'b1;
 		default: edge_mask_reg_p6[97] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110011,
	14'b1001011110100,
	14'b1001011110101,
	14'b1001100000011,
	14'b1001100000100,
	14'b1001100000101,
	14'b1001100010011,
	14'b1001100010100,
	14'b1001100010101,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100010101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100010101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10001011100000,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10101100000000: edge_mask_reg_p6[98] <= 1'b1;
 		default: edge_mask_reg_p6[98] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110100,
	14'b1001011110101,
	14'b1001011110110,
	14'b1001100000100,
	14'b1001100000101,
	14'b1001100000110,
	14'b1001100010100,
	14'b1001100010101,
	14'b1001100010110,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100010110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100010110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10001011100000,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[99] <= 1'b1;
 		default: edge_mask_reg_p6[99] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110101,
	14'b1001011110110,
	14'b1001011110111,
	14'b1001100000101,
	14'b1001100000110,
	14'b1001100000111,
	14'b1001100010101,
	14'b1001100010110,
	14'b1001100010111,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100010101,
	14'b1010100010110,
	14'b1010100010111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100010111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[100] <= 1'b1;
 		default: edge_mask_reg_p6[100] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001011110110,
	14'b1001011110111,
	14'b1001011111000,
	14'b1001100000110,
	14'b1001100000111,
	14'b1001100001000,
	14'b1001100010110,
	14'b1001100010111,
	14'b1001100011000,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010011111000,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100001000,
	14'b1010100010110,
	14'b1010100010111,
	14'b1010100011000,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100011000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110000,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000: edge_mask_reg_p6[101] <= 1'b1;
 		default: edge_mask_reg_p6[101] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110111,
	14'b1010011111000,
	14'b1010011111001,
	14'b1010100000111,
	14'b1010100001000,
	14'b1010100001001,
	14'b1010100010111,
	14'b1010100011000,
	14'b1010100011001,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100011001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1110011100000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[102] <= 1'b1;
 		default: edge_mask_reg_p6[102] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011111000,
	14'b1010011111001,
	14'b1010011111010,
	14'b1010100001000,
	14'b1010100001001,
	14'b1010100001010,
	14'b1010100011000,
	14'b1010100011001,
	14'b1010100011010,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101011111011,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100001011,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100011011,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100001011,
	14'b1110100010000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101100000001,
	14'b10101100010001: edge_mask_reg_p6[103] <= 1'b1;
 		default: edge_mask_reg_p6[103] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100010000,
	14'b1001100100000,
	14'b1001100110000,
	14'b1010100010000,
	14'b1010100100000,
	14'b1010100110000,
	14'b1011100010000,
	14'b1011100100000,
	14'b1011100110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100110000: edge_mask_reg_p6[104] <= 1'b1;
 		default: edge_mask_reg_p6[104] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100010000,
	14'b1001100010001,
	14'b1001100100000,
	14'b1001100100001,
	14'b1001100110000,
	14'b1001100110001,
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100110000,
	14'b1010100110001,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10001011110000,
	14'b10001100000000: edge_mask_reg_p6[105] <= 1'b1;
 		default: edge_mask_reg_p6[105] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100010000,
	14'b1001100010001,
	14'b1001100010010,
	14'b1001100100000,
	14'b1001100100001,
	14'b1001100100010,
	14'b1001100110000,
	14'b1001100110001,
	14'b1001100110010,
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10010011110000,
	14'b10010100000000: edge_mask_reg_p6[106] <= 1'b1;
 		default: edge_mask_reg_p6[106] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000001,
	14'b1001100000010,
	14'b1001100000011,
	14'b1001100010001,
	14'b1001100010010,
	14'b1001100010011,
	14'b1001100100001,
	14'b1001100100010,
	14'b1001100100011,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[107] <= 1'b1;
 		default: edge_mask_reg_p6[107] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000010,
	14'b1001100000011,
	14'b1001100000100,
	14'b1001100010010,
	14'b1001100010011,
	14'b1001100010100,
	14'b1001100100010,
	14'b1001100100011,
	14'b1001100100100,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100100100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000010,
	14'b10000101000011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011100000000,
	14'b10011100010000: edge_mask_reg_p6[108] <= 1'b1;
 		default: edge_mask_reg_p6[108] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000011,
	14'b1001100000100,
	14'b1001100000101,
	14'b1001100010011,
	14'b1001100010100,
	14'b1001100010101,
	14'b1001100100011,
	14'b1001100100100,
	14'b1001100100101,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100100101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100100101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000011,
	14'b10000101000100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[109] <= 1'b1;
 		default: edge_mask_reg_p6[109] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000100,
	14'b1001100000101,
	14'b1001100000110,
	14'b1001100010100,
	14'b1001100010101,
	14'b1001100010110,
	14'b1001100100100,
	14'b1001100100101,
	14'b1001100100110,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100010110,
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100100110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100100110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000100,
	14'b10000101000101,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110010,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[110] <= 1'b1;
 		default: edge_mask_reg_p6[110] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000101,
	14'b1001100000110,
	14'b1001100000111,
	14'b1001100010101,
	14'b1001100010110,
	14'b1001100010111,
	14'b1001100100101,
	14'b1001100100110,
	14'b1001100100111,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100010101,
	14'b1010100010110,
	14'b1010100010111,
	14'b1010100100101,
	14'b1010100100110,
	14'b1010100100111,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100100111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[111] <= 1'b1;
 		default: edge_mask_reg_p6[111] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100000110,
	14'b1001100000111,
	14'b1001100001000,
	14'b1001100010110,
	14'b1001100010111,
	14'b1001100011000,
	14'b1001100100110,
	14'b1001100100111,
	14'b1001100101000,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100001000,
	14'b1010100010110,
	14'b1010100010111,
	14'b1010100011000,
	14'b1010100100110,
	14'b1010100100111,
	14'b1010100101000,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100101000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000: edge_mask_reg_p6[112] <= 1'b1;
 		default: edge_mask_reg_p6[112] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100000111,
	14'b1010100001000,
	14'b1010100001001,
	14'b1010100010111,
	14'b1010100011000,
	14'b1010100011001,
	14'b1010100100111,
	14'b1010100101000,
	14'b1010100101001,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100101001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[113] <= 1'b1;
 		default: edge_mask_reg_p6[113] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100001000,
	14'b1010100001001,
	14'b1010100001010,
	14'b1010100011000,
	14'b1010100011001,
	14'b1010100011010,
	14'b1010100101000,
	14'b1010100101001,
	14'b1010100101010,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100101010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100011011,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100101011,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110000,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[114] <= 1'b1;
 		default: edge_mask_reg_p6[114] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100000,
	14'b1001100110000,
	14'b1001101000000,
	14'b1010100100000,
	14'b1010100110000,
	14'b1010101000000,
	14'b1011100100000,
	14'b1011100110000,
	14'b1011101000000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000: edge_mask_reg_p6[115] <= 1'b1;
 		default: edge_mask_reg_p6[115] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100000,
	14'b1001100100001,
	14'b1001100110000,
	14'b1001100110001,
	14'b1001101000000,
	14'b1001101000001,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010101000000,
	14'b1010101000001,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100000000,
	14'b10001100010000: edge_mask_reg_p6[116] <= 1'b1;
 		default: edge_mask_reg_p6[116] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100000,
	14'b1001100100001,
	14'b1001100100010,
	14'b1001100110000,
	14'b1001100110001,
	14'b1001100110010,
	14'b1001101000000,
	14'b1001101000001,
	14'b1001101000010,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10010100000000,
	14'b10010100010000: edge_mask_reg_p6[117] <= 1'b1;
 		default: edge_mask_reg_p6[117] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100001,
	14'b1001100100010,
	14'b1001100100011,
	14'b1001100110001,
	14'b1001100110010,
	14'b1001100110011,
	14'b1001101000001,
	14'b1001101000010,
	14'b1001101000011,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010001,
	14'b1111101010010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010001,
	14'b10000101010010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[118] <= 1'b1;
 		default: edge_mask_reg_p6[118] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100010,
	14'b1001100100011,
	14'b1001100100100,
	14'b1001100110010,
	14'b1001100110011,
	14'b1001100110100,
	14'b1001101000010,
	14'b1001101000011,
	14'b1001101000100,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010010,
	14'b10000101010011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[119] <= 1'b1;
 		default: edge_mask_reg_p6[119] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100011,
	14'b1001100100100,
	14'b1001100100101,
	14'b1001100110011,
	14'b1001100110100,
	14'b1001100110101,
	14'b1001101000011,
	14'b1001101000100,
	14'b1001101000101,
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010011,
	14'b10000101010100,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[120] <= 1'b1;
 		default: edge_mask_reg_p6[120] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100100,
	14'b1001100100101,
	14'b1001100100110,
	14'b1001100110100,
	14'b1001100110101,
	14'b1001100110110,
	14'b1001101000100,
	14'b1001101000101,
	14'b1001101000110,
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100100110,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010100110110,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101000110,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010100,
	14'b10000101010101,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[121] <= 1'b1;
 		default: edge_mask_reg_p6[121] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100101,
	14'b1001100100110,
	14'b1001100100111,
	14'b1001100110101,
	14'b1001100110110,
	14'b1001100110111,
	14'b1001101000101,
	14'b1001101000110,
	14'b1001101000111,
	14'b1010100100101,
	14'b1010100100110,
	14'b1010100100111,
	14'b1010100110101,
	14'b1010100110110,
	14'b1010100110111,
	14'b1010101000101,
	14'b1010101000110,
	14'b1010101000111,
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010101,
	14'b10000101010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[122] <= 1'b1;
 		default: edge_mask_reg_p6[122] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100100110,
	14'b1001100100111,
	14'b1001100101000,
	14'b1001100110110,
	14'b1001100110111,
	14'b1001100111000,
	14'b1001101000110,
	14'b1001101000111,
	14'b1001101001000,
	14'b1010100100110,
	14'b1010100100111,
	14'b1010100101000,
	14'b1010100110110,
	14'b1010100110111,
	14'b1010100111000,
	14'b1010101000110,
	14'b1010101000111,
	14'b1010101001000,
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010110,
	14'b10000101010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[123] <= 1'b1;
 		default: edge_mask_reg_p6[123] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100111,
	14'b1010100101000,
	14'b1010100101001,
	14'b1010100110111,
	14'b1010100111000,
	14'b1010100111001,
	14'b1010101000111,
	14'b1010101001000,
	14'b1010101001001,
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100001: edge_mask_reg_p6[124] <= 1'b1;
 		default: edge_mask_reg_p6[124] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100011000,
	14'b1010100011001,
	14'b1010100011010,
	14'b1010100101000,
	14'b1010100101001,
	14'b1010100101010,
	14'b1010100111000,
	14'b1010100111001,
	14'b1010100111010,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100101010,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011100111010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100011011,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100101011,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101100111011,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010: edge_mask_reg_p6[125] <= 1'b1;
 		default: edge_mask_reg_p6[125] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110000,
	14'b1001101000000,
	14'b1001101010000,
	14'b1010100110000,
	14'b1010101000000,
	14'b1010101010000,
	14'b1011100110000,
	14'b1011101000000,
	14'b1011101010000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1100101010000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1110100010000,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100100000: edge_mask_reg_p6[126] <= 1'b1;
 		default: edge_mask_reg_p6[126] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110000,
	14'b1001100110001,
	14'b1001101000000,
	14'b1001101000001,
	14'b1001101010000,
	14'b1001101010001,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101010000,
	14'b1010101010001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100010000,
	14'b10001100100000: edge_mask_reg_p6[127] <= 1'b1;
 		default: edge_mask_reg_p6[127] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110000,
	14'b1001100110001,
	14'b1001100110010,
	14'b1001101000000,
	14'b1001101000001,
	14'b1001101000010,
	14'b1001101010000,
	14'b1001101010001,
	14'b1001101010010,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101010000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[128] <= 1'b1;
 		default: edge_mask_reg_p6[128] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110001,
	14'b1001100110010,
	14'b1001100110011,
	14'b1001101000001,
	14'b1001101000010,
	14'b1001101000011,
	14'b1001101010001,
	14'b1001101010010,
	14'b1001101010011,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100001,
	14'b1111101100010,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100001,
	14'b10000101100010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010101000000: edge_mask_reg_p6[129] <= 1'b1;
 		default: edge_mask_reg_p6[129] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110010,
	14'b1001100110011,
	14'b1001100110100,
	14'b1001101000010,
	14'b1001101000011,
	14'b1001101000100,
	14'b1001101010010,
	14'b1001101010011,
	14'b1001101010100,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100010,
	14'b1111101100011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100010,
	14'b10000101100011,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010001,
	14'b10001101010010,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011110000: edge_mask_reg_p6[130] <= 1'b1;
 		default: edge_mask_reg_p6[130] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110011,
	14'b1001100110100,
	14'b1001100110101,
	14'b1001101000011,
	14'b1001101000100,
	14'b1001101000101,
	14'b1001101010011,
	14'b1001101010100,
	14'b1001101010101,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100011,
	14'b1111101100100,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100011,
	14'b10000101100100,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010010,
	14'b10001101010011,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[131] <= 1'b1;
 		default: edge_mask_reg_p6[131] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110100,
	14'b1001100110101,
	14'b1001100110110,
	14'b1001101000100,
	14'b1001101000101,
	14'b1001101000110,
	14'b1001101010100,
	14'b1001101010101,
	14'b1001101010110,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010100110110,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101000110,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101010110,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100100,
	14'b10000101100101,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010011,
	14'b10001101010100,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[132] <= 1'b1;
 		default: edge_mask_reg_p6[132] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110101,
	14'b1001100110110,
	14'b1001100110111,
	14'b1001101000101,
	14'b1001101000110,
	14'b1001101000111,
	14'b1001101010101,
	14'b1001101010110,
	14'b1001101010111,
	14'b1010100110101,
	14'b1010100110110,
	14'b1010100110111,
	14'b1010101000101,
	14'b1010101000110,
	14'b1010101000111,
	14'b1010101010101,
	14'b1010101010110,
	14'b1010101010111,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100101,
	14'b10000101100110,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000010,
	14'b10010101000011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[133] <= 1'b1;
 		default: edge_mask_reg_p6[133] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001100110110,
	14'b1001100110111,
	14'b1001100111000,
	14'b1001101000110,
	14'b1001101000111,
	14'b1001101001000,
	14'b1001101010110,
	14'b1001101010111,
	14'b1001101011000,
	14'b1010100110110,
	14'b1010100110111,
	14'b1010100111000,
	14'b1010101000110,
	14'b1010101000111,
	14'b1010101001000,
	14'b1010101010110,
	14'b1010101010111,
	14'b1010101011000,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1110011110000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100110,
	14'b10000101100111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000011,
	14'b10010101000100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[134] <= 1'b1;
 		default: edge_mask_reg_p6[134] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110111,
	14'b1010100111000,
	14'b1010100111001,
	14'b1010101000111,
	14'b1010101001000,
	14'b1010101001001,
	14'b1010101010111,
	14'b1010101011000,
	14'b1010101011001,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100111,
	14'b10000101101000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[135] <= 1'b1;
 		default: edge_mask_reg_p6[135] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100111000,
	14'b1010100111001,
	14'b1010100111010,
	14'b1010101001000,
	14'b1010101001001,
	14'b1010101001010,
	14'b1010101011000,
	14'b1010101011001,
	14'b1010101011010,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011100111010,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101001010,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100101011,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101100111011,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101001011,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101101000,
	14'b10000101101001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010110,
	14'b10001101010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010: edge_mask_reg_p6[136] <= 1'b1;
 		default: edge_mask_reg_p6[136] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000000,
	14'b1001101010000,
	14'b1001101100000,
	14'b1010101000000,
	14'b1010101010000,
	14'b1010101100000,
	14'b1011101000000,
	14'b1011101010000,
	14'b1011101100000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101100000,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101100000,
	14'b10001100100000,
	14'b10001100110000: edge_mask_reg_p6[137] <= 1'b1;
 		default: edge_mask_reg_p6[137] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000000,
	14'b1001101000001,
	14'b1001101010000,
	14'b1001101010001,
	14'b1001101100000,
	14'b1001101100001,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101100000,
	14'b1010101100001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010100100000: edge_mask_reg_p6[138] <= 1'b1;
 		default: edge_mask_reg_p6[138] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000000,
	14'b1001101000001,
	14'b1001101000010,
	14'b1001101010000,
	14'b1001101010001,
	14'b1001101010010,
	14'b1001101100000,
	14'b1001101100001,
	14'b1001101100010,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101010000,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[139] <= 1'b1;
 		default: edge_mask_reg_p6[139] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000001,
	14'b1001101000010,
	14'b1001101000011,
	14'b1001101010001,
	14'b1001101010010,
	14'b1001101010011,
	14'b1001101100001,
	14'b1001101100010,
	14'b1001101100011,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110001,
	14'b1111101110010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110001,
	14'b10000101110010,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000: edge_mask_reg_p6[140] <= 1'b1;
 		default: edge_mask_reg_p6[140] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000010,
	14'b1001101000011,
	14'b1001101000100,
	14'b1001101010010,
	14'b1001101010011,
	14'b1001101010100,
	14'b1001101100010,
	14'b1001101100011,
	14'b1001101100100,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110010,
	14'b1111101110011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110010,
	14'b10000101110011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100001,
	14'b10001101100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[141] <= 1'b1;
 		default: edge_mask_reg_p6[141] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000011,
	14'b1001101000100,
	14'b1001101000101,
	14'b1001101010011,
	14'b1001101010100,
	14'b1001101010101,
	14'b1001101100011,
	14'b1001101100100,
	14'b1001101100101,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101100101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110011,
	14'b1111101110100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110011,
	14'b10000101110100,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100010,
	14'b10001101100011,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[142] <= 1'b1;
 		default: edge_mask_reg_p6[142] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000100,
	14'b1001101000101,
	14'b1001101000110,
	14'b1001101010100,
	14'b1001101010101,
	14'b1001101010110,
	14'b1001101100100,
	14'b1001101100101,
	14'b1001101100110,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101000110,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101010110,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101100110,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1100100110101,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110100,
	14'b1111101110101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110100,
	14'b10000101110101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100011,
	14'b10001101100100,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000: edge_mask_reg_p6[143] <= 1'b1;
 		default: edge_mask_reg_p6[143] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101000101,
	14'b1001101000110,
	14'b1001101000111,
	14'b1001101010101,
	14'b1001101010110,
	14'b1001101010111,
	14'b1001101100101,
	14'b1001101100110,
	14'b1001101100111,
	14'b1010101000101,
	14'b1010101000110,
	14'b1010101000111,
	14'b1010101010101,
	14'b1010101010110,
	14'b1010101010111,
	14'b1010101100101,
	14'b1010101100110,
	14'b1010101100111,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1100100110110,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110101,
	14'b1111101110110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110101,
	14'b10000101110110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[144] <= 1'b1;
 		default: edge_mask_reg_p6[144] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000110,
	14'b1010101000111,
	14'b1010101001000,
	14'b1010101010110,
	14'b1010101010111,
	14'b1010101011000,
	14'b1010101100110,
	14'b1010101100111,
	14'b1010101101000,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110110,
	14'b10000101110111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[145] <= 1'b1;
 		default: edge_mask_reg_p6[145] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000111,
	14'b1010101001000,
	14'b1010101001001,
	14'b1010101010111,
	14'b1010101011000,
	14'b1010101011001,
	14'b1010101100111,
	14'b1010101101000,
	14'b1010101101001,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1101011110000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110111,
	14'b10000101111000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[146] <= 1'b1;
 		default: edge_mask_reg_p6[146] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101001000,
	14'b1010101001001,
	14'b1010101001010,
	14'b1010101011000,
	14'b1010101011001,
	14'b1010101011010,
	14'b1010101101000,
	14'b1010101101001,
	14'b1010101101010,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101001010,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101100111011,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101001011,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101011011,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000000,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101111000,
	14'b10000101111001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110010: edge_mask_reg_p6[147] <= 1'b1;
 		default: edge_mask_reg_p6[147] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010000,
	14'b1001101100000,
	14'b1001101110000,
	14'b1010101010000,
	14'b1010101100000,
	14'b1010101110000,
	14'b1011101010000,
	14'b1011101100000,
	14'b1011101110000,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101110000,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101010000: edge_mask_reg_p6[148] <= 1'b1;
 		default: edge_mask_reg_p6[148] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010000,
	14'b1001101010001,
	14'b1001101100000,
	14'b1001101100001,
	14'b1001101110000,
	14'b1001101110001,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101110000,
	14'b1010101110001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010100110000: edge_mask_reg_p6[149] <= 1'b1;
 		default: edge_mask_reg_p6[149] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010000,
	14'b1001101010001,
	14'b1001101010010,
	14'b1001101100000,
	14'b1001101100001,
	14'b1001101100010,
	14'b1001101110000,
	14'b1001101110001,
	14'b1001101110010,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101100000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000: edge_mask_reg_p6[150] <= 1'b1;
 		default: edge_mask_reg_p6[150] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010001,
	14'b1001101010010,
	14'b1001101010011,
	14'b1001101100001,
	14'b1001101100010,
	14'b1001101100011,
	14'b1001101110001,
	14'b1001101110010,
	14'b1001101110011,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000001,
	14'b1111110000010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10010100000000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101100000000: edge_mask_reg_p6[151] <= 1'b1;
 		default: edge_mask_reg_p6[151] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010010,
	14'b1001101010011,
	14'b1001101010100,
	14'b1001101100010,
	14'b1001101100011,
	14'b1001101100100,
	14'b1001101110010,
	14'b1001101110011,
	14'b1001101110100,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010101110100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000010,
	14'b1111110000011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000010,
	14'b10000110000011,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[152] <= 1'b1;
 		default: edge_mask_reg_p6[152] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010011,
	14'b1001101010100,
	14'b1001101010101,
	14'b1001101100011,
	14'b1001101100100,
	14'b1001101100101,
	14'b1001101110011,
	14'b1001101110100,
	14'b1001101110101,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010101110101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000011,
	14'b1111110000100,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000011,
	14'b10000110000100,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[153] <= 1'b1;
 		default: edge_mask_reg_p6[153] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010100,
	14'b1001101010101,
	14'b1001101010110,
	14'b1001101100100,
	14'b1001101100101,
	14'b1001101100110,
	14'b1001101110100,
	14'b1001101110101,
	14'b1001101110110,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101010110,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101100110,
	14'b1010101110100,
	14'b1010101110101,
	14'b1010101110110,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1100101000101,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000100,
	14'b1111110000101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000100,
	14'b10000110000101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[154] <= 1'b1;
 		default: edge_mask_reg_p6[154] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101010101,
	14'b1001101010110,
	14'b1001101010111,
	14'b1001101100101,
	14'b1001101100110,
	14'b1001101100111,
	14'b1001101110101,
	14'b1001101110110,
	14'b1001101110111,
	14'b1010101010101,
	14'b1010101010110,
	14'b1010101010111,
	14'b1010101100101,
	14'b1010101100110,
	14'b1010101100111,
	14'b1010101110101,
	14'b1010101110110,
	14'b1010101110111,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1100101000110,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100100100,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000101,
	14'b1111110000110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000101,
	14'b10000110000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[155] <= 1'b1;
 		default: edge_mask_reg_p6[155] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010110,
	14'b1010101010111,
	14'b1010101011000,
	14'b1010101100110,
	14'b1010101100111,
	14'b1010101101000,
	14'b1010101110110,
	14'b1010101110111,
	14'b1010101111000,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1100101000111,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000110,
	14'b1111110000111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000110,
	14'b10000110000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000: edge_mask_reg_p6[156] <= 1'b1;
 		default: edge_mask_reg_p6[156] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010111,
	14'b1010101011000,
	14'b1010101011001,
	14'b1010101100111,
	14'b1010101101000,
	14'b1010101101001,
	14'b1010101110111,
	14'b1010101111000,
	14'b1010101111001,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000111,
	14'b1111110001000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000111,
	14'b10000110001000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[157] <= 1'b1;
 		default: edge_mask_reg_p6[157] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101011000,
	14'b1010101011001,
	14'b1010101011010,
	14'b1010101101000,
	14'b1010101101001,
	14'b1010101101010,
	14'b1010101111000,
	14'b1010101111001,
	14'b1010101111010,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1100011110000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101001011,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101011011,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101101011,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100110,
	14'b1110100110000,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010000,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110001000,
	14'b10000110001001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[158] <= 1'b1;
 		default: edge_mask_reg_p6[158] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100000,
	14'b1001101110000,
	14'b1001110000000,
	14'b1010101100000,
	14'b1010101110000,
	14'b1010110000000,
	14'b1011101100000,
	14'b1011101110000,
	14'b1011110000000,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100110000000,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101100000: edge_mask_reg_p6[159] <= 1'b1;
 		default: edge_mask_reg_p6[159] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100000,
	14'b1001101100001,
	14'b1001101110000,
	14'b1001101110001,
	14'b1001110000000,
	14'b1001110000001,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010110000000,
	14'b1010110000001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011110000000,
	14'b1011110000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100001,
	14'b10010100110000,
	14'b10010101000000: edge_mask_reg_p6[160] <= 1'b1;
 		default: edge_mask_reg_p6[160] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100000,
	14'b1001101100001,
	14'b1001101100010,
	14'b1001101110000,
	14'b1001101110001,
	14'b1001101110010,
	14'b1001110000000,
	14'b1001110000001,
	14'b1001110000010,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110000010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110000010,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110010000,
	14'b1101110010001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101110000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011100010000,
	14'b10100100010000: edge_mask_reg_p6[161] <= 1'b1;
 		default: edge_mask_reg_p6[161] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100001,
	14'b1001101100010,
	14'b1001101100011,
	14'b1001101110001,
	14'b1001101110010,
	14'b1001101110011,
	14'b1001110000001,
	14'b1001110000010,
	14'b1001110000011,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110000011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110000011,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110010001,
	14'b1101110010010,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010001,
	14'b1110110010010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[162] <= 1'b1;
 		default: edge_mask_reg_p6[162] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100010,
	14'b1001101100011,
	14'b1001101100100,
	14'b1001101110010,
	14'b1001101110011,
	14'b1001101110100,
	14'b1001110000010,
	14'b1001110000011,
	14'b1001110000100,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010110000010,
	14'b1010110000011,
	14'b1010110000100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110000100,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110010010,
	14'b1101110010011,
	14'b1110100110010,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010010,
	14'b1110110010011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010010,
	14'b1111110010011,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010010,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[163] <= 1'b1;
 		default: edge_mask_reg_p6[163] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100011,
	14'b1001101100100,
	14'b1001101100101,
	14'b1001101110011,
	14'b1001101110100,
	14'b1001101110101,
	14'b1001110000011,
	14'b1001110000100,
	14'b1001110000101,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010101110101,
	14'b1010110000011,
	14'b1010110000100,
	14'b1010110000101,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110000101,
	14'b1100101010100,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110010011,
	14'b1101110010100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010011,
	14'b1110110010100,
	14'b1111100000000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010011,
	14'b1111110010100,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010011,
	14'b10000110010100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[164] <= 1'b1;
 		default: edge_mask_reg_p6[164] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101100100,
	14'b1001101100101,
	14'b1001101100110,
	14'b1001101110100,
	14'b1001101110101,
	14'b1001101110110,
	14'b1001110000100,
	14'b1001110000101,
	14'b1001110000110,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101100110,
	14'b1010101110100,
	14'b1010101110101,
	14'b1010101110110,
	14'b1010110000100,
	14'b1010110000101,
	14'b1010110000110,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110000110,
	14'b1100101010101,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110010100,
	14'b1101110010101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010100,
	14'b1110110010101,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010100,
	14'b1111110010101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010100,
	14'b10000110010101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100001,
	14'b10010101100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[165] <= 1'b1;
 		default: edge_mask_reg_p6[165] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100101,
	14'b1010101100110,
	14'b1010101100111,
	14'b1010101110101,
	14'b1010101110110,
	14'b1010101110111,
	14'b1010110000101,
	14'b1010110000110,
	14'b1010110000111,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110000111,
	14'b1100101010110,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110010101,
	14'b1101110010110,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010101,
	14'b1110110010110,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010101,
	14'b1111110010110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010101,
	14'b10000110010110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110011,
	14'b10001101110100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100010,
	14'b10010101100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101100110001,
	14'b10101101000000: edge_mask_reg_p6[166] <= 1'b1;
 		default: edge_mask_reg_p6[166] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100110,
	14'b1010101100111,
	14'b1010101101000,
	14'b1010101110110,
	14'b1010101110111,
	14'b1010101111000,
	14'b1010110000110,
	14'b1010110000111,
	14'b1010110001000,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110001000,
	14'b1100101010111,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1101100000000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110010110,
	14'b1101110010111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010110,
	14'b1110110010111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010110,
	14'b1111110010111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010110,
	14'b10000110010111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[167] <= 1'b1;
 		default: edge_mask_reg_p6[167] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100111,
	14'b1010101101000,
	14'b1010101101001,
	14'b1010101110111,
	14'b1010101111000,
	14'b1010101111001,
	14'b1010110000111,
	14'b1010110001000,
	14'b1010110001001,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110001001,
	14'b1100101011000,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110010111,
	14'b1101110011000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010111,
	14'b1110110011000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010111,
	14'b1111110011000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010111,
	14'b10000110011000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000001,
	14'b10100101000010: edge_mask_reg_p6[168] <= 1'b1;
 		default: edge_mask_reg_p6[168] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101101000,
	14'b1010101101001,
	14'b1010101101010,
	14'b1010101111000,
	14'b1010101111001,
	14'b1010101111010,
	14'b1010110001000,
	14'b1010110001001,
	14'b1010110001010,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110001010,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100101011001,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101101000000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101011011,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101101011,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101101111011,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110011000,
	14'b1101110011001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110101111011,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110011000,
	14'b1110110011001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110011000,
	14'b1111110011001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110011000,
	14'b10000110011001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110101,
	14'b10001101110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100001,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011: edge_mask_reg_p6[169] <= 1'b1;
 		default: edge_mask_reg_p6[169] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110000,
	14'b1001110000000,
	14'b1001110010000,
	14'b1010101110000,
	14'b1010110000000,
	14'b1010110010000,
	14'b1011101110000,
	14'b1011110000000,
	14'b1011110010000,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110010000,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110010000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111101010000,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000101010000,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110010000,
	14'b10001101010000,
	14'b10001101100000,
	14'b10001101110000: edge_mask_reg_p6[170] <= 1'b1;
 		default: edge_mask_reg_p6[170] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110000,
	14'b1001101110001,
	14'b1001110000000,
	14'b1001110000001,
	14'b1001110010000,
	14'b1001110010001,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110010000,
	14'b1010110010001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110010000,
	14'b1011110010001,
	14'b1100101100000,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110010000,
	14'b1100110010001,
	14'b1101101010000,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110010000,
	14'b1101110010001,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110001,
	14'b10010101000000,
	14'b10010101010000: edge_mask_reg_p6[171] <= 1'b1;
 		default: edge_mask_reg_p6[171] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110000,
	14'b1001101110001,
	14'b1001101110010,
	14'b1001110000000,
	14'b1001110000001,
	14'b1001110000010,
	14'b1001110010000,
	14'b1001110010001,
	14'b1001110010010,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110010000,
	14'b1010110010001,
	14'b1010110010010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110010000,
	14'b1011110010001,
	14'b1011110010010,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110010000,
	14'b1100110010001,
	14'b1100110010010,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110010000,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110100000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110100000,
	14'b1110110100001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110100000,
	14'b1111110100001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001110000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[172] <= 1'b1;
 		default: edge_mask_reg_p6[172] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110001,
	14'b1001101110010,
	14'b1001101110011,
	14'b1001110000001,
	14'b1001110000010,
	14'b1001110000011,
	14'b1001110010001,
	14'b1001110010010,
	14'b1001110010011,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110000011,
	14'b1010110010001,
	14'b1010110010010,
	14'b1010110010011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110010001,
	14'b1011110010010,
	14'b1011110010011,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110010001,
	14'b1100110010010,
	14'b1100110010011,
	14'b1101101010010,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110010000,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110100001,
	14'b1101110100010,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110100001,
	14'b1110110100010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110100001,
	14'b1111110100010,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110100001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[173] <= 1'b1;
 		default: edge_mask_reg_p6[173] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110010,
	14'b1001101110011,
	14'b1001101110100,
	14'b1001110000010,
	14'b1001110000011,
	14'b1001110000100,
	14'b1001110010010,
	14'b1001110010011,
	14'b1001110010100,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010110000010,
	14'b1010110000011,
	14'b1010110000100,
	14'b1010110010010,
	14'b1010110010011,
	14'b1010110010100,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110010010,
	14'b1011110010011,
	14'b1011110010100,
	14'b1100101100011,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110010010,
	14'b1100110010011,
	14'b1100110010100,
	14'b1101101010011,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110100010,
	14'b1101110100011,
	14'b1110101000010,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110100010,
	14'b1110110100011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110100010,
	14'b1111110100011,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110100010,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101010000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[174] <= 1'b1;
 		default: edge_mask_reg_p6[174] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1001101110011,
	14'b1001101110100,
	14'b1001101110101,
	14'b1001110000011,
	14'b1001110000100,
	14'b1001110000101,
	14'b1001110010011,
	14'b1001110010100,
	14'b1001110010101,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010101110101,
	14'b1010110000011,
	14'b1010110000100,
	14'b1010110000101,
	14'b1010110010011,
	14'b1010110010100,
	14'b1010110010101,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110010011,
	14'b1011110010100,
	14'b1011110010101,
	14'b1100101100100,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110010011,
	14'b1100110010100,
	14'b1100110010101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110100011,
	14'b1101110100100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110100011,
	14'b1110110100100,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110100011,
	14'b1111110100100,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110100011,
	14'b10000110100100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000001,
	14'b10001110000010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[175] <= 1'b1;
 		default: edge_mask_reg_p6[175] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110100,
	14'b1010101110101,
	14'b1010101110110,
	14'b1010110000100,
	14'b1010110000101,
	14'b1010110000110,
	14'b1010110010100,
	14'b1010110010101,
	14'b1010110010110,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110010100,
	14'b1011110010101,
	14'b1011110010110,
	14'b1100101100101,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110010100,
	14'b1100110010101,
	14'b1100110010110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110100100,
	14'b1101110100101,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110100100,
	14'b1110110100101,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110100100,
	14'b1111110100101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110100100,
	14'b10000110100101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000010,
	14'b10001110000011,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110001,
	14'b10010101110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[176] <= 1'b1;
 		default: edge_mask_reg_p6[176] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110101,
	14'b1010101110110,
	14'b1010101110111,
	14'b1010110000101,
	14'b1010110000110,
	14'b1010110000111,
	14'b1010110010101,
	14'b1010110010110,
	14'b1010110010111,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110010101,
	14'b1011110010110,
	14'b1011110010111,
	14'b1100101100110,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110010101,
	14'b1100110010110,
	14'b1100110010111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110100101,
	14'b1101110100110,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110100101,
	14'b1110110100110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110100101,
	14'b1111110100110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110100101,
	14'b10000110100110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000011,
	14'b10001110000100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10100101010001,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[177] <= 1'b1;
 		default: edge_mask_reg_p6[177] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110110,
	14'b1010101110111,
	14'b1010101111000,
	14'b1010110000110,
	14'b1010110000111,
	14'b1010110001000,
	14'b1010110010110,
	14'b1010110010111,
	14'b1010110011000,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110010110,
	14'b1011110010111,
	14'b1011110011000,
	14'b1100101100111,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110010110,
	14'b1100110010111,
	14'b1100110011000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110100110,
	14'b1101110100111,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110100110,
	14'b1110110100111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110100110,
	14'b1111110100111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110100110,
	14'b10000110100111,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000100,
	14'b10001110000101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010: edge_mask_reg_p6[178] <= 1'b1;
 		default: edge_mask_reg_p6[178] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110111,
	14'b1010101111000,
	14'b1010101111001,
	14'b1010110000111,
	14'b1010110001000,
	14'b1010110001001,
	14'b1010110010111,
	14'b1010110011000,
	14'b1010110011001,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110010111,
	14'b1011110011000,
	14'b1011110011001,
	14'b1100100000000,
	14'b1100101101000,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110010111,
	14'b1100110011000,
	14'b1100110011001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110011001,
	14'b1101110100111,
	14'b1101110101000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010000,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110100111,
	14'b1110110101000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110100111,
	14'b1111110101000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110100111,
	14'b10000110101000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000: edge_mask_reg_p6[179] <= 1'b1;
 		default: edge_mask_reg_p6[179] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101111000,
	14'b1010101111001,
	14'b1010101111010,
	14'b1010110001000,
	14'b1010110001001,
	14'b1010110001010,
	14'b1010110011000,
	14'b1010110011001,
	14'b1010110011010,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110001010,
	14'b1011110011000,
	14'b1011110011001,
	14'b1011110011010,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100101101001,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1100110011000,
	14'b1100110011001,
	14'b1100110011010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100010,
	14'b1101101000000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010000,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101101011,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101101111011,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110001011,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110011001,
	14'b1101110011010,
	14'b1101110101000,
	14'b1101110101001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110101111011,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110001011,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110011010,
	14'b1110110101000,
	14'b1110110101001,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110001011,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110011010,
	14'b1111110101000,
	14'b1111110101001,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110001011,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110011010,
	14'b10000110101000,
	14'b10000110101001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010100000010,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010: edge_mask_reg_p6[180] <= 1'b1;
 		default: edge_mask_reg_p6[180] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100000,
	14'b1010001110000,
	14'b1010010000000,
	14'b1011001100000,
	14'b1011001110000,
	14'b1011010000000,
	14'b1100001100000,
	14'b1100001110000,
	14'b1100010000000,
	14'b1101001100000,
	14'b1101001110000,
	14'b1101010000000,
	14'b1110001100000,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10010010010000,
	14'b10010010100000: edge_mask_reg_p6[181] <= 1'b1;
 		default: edge_mask_reg_p6[181] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100000,
	14'b1010001100001,
	14'b1010001110000,
	14'b1010001110001,
	14'b1010010000000,
	14'b1010010000001,
	14'b1011001100000,
	14'b1011001100001,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011010000000,
	14'b1011010000001,
	14'b1100001100000,
	14'b1100001100001,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1110001010000,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1111001010000,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b10000001010000,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010110000: edge_mask_reg_p6[182] <= 1'b1;
 		default: edge_mask_reg_p6[182] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100000,
	14'b1010001100001,
	14'b1010001100010,
	14'b1010001110000,
	14'b1010001110001,
	14'b1010001110010,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010000010,
	14'b1011001100000,
	14'b1011001100001,
	14'b1011001100010,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010000010,
	14'b1100001100000,
	14'b1100001100001,
	14'b1100001100010,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1110001010000,
	14'b1110001010001,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1111001010000,
	14'b1111001010001,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b10000001010000,
	14'b10000001010001,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10001001010000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10010010000000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10011010100000,
	14'b10011010110000: edge_mask_reg_p6[183] <= 1'b1;
 		default: edge_mask_reg_p6[183] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001100001,
	14'b1010001100010,
	14'b1010001100011,
	14'b1010001110001,
	14'b1010001110010,
	14'b1010001110011,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010000011,
	14'b1011001100001,
	14'b1011001100010,
	14'b1011001100011,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010000011,
	14'b1100001100001,
	14'b1100001100010,
	14'b1100001100011,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1110001010001,
	14'b1110001010010,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100001,
	14'b1110010100010,
	14'b1111001010001,
	14'b1111001010010,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b10000001010001,
	14'b10000001010010,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001001010001,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001110000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10101011100000: edge_mask_reg_p6[184] <= 1'b1;
 		default: edge_mask_reg_p6[184] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100010,
	14'b1011001100011,
	14'b1011001100100,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011001110100,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010000100,
	14'b1100001100010,
	14'b1100001100011,
	14'b1100001100100,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1110001010010,
	14'b1110001010011,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100010,
	14'b1110010100011,
	14'b1111001010010,
	14'b1111001010011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110001,
	14'b1111010110010,
	14'b10000001010010,
	14'b10000001010011,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10001001010010,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10101011010000,
	14'b10101011100000: edge_mask_reg_p6[185] <= 1'b1;
 		default: edge_mask_reg_p6[185] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100011,
	14'b1011001100100,
	14'b1011001100101,
	14'b1011001110011,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010000101,
	14'b1100001100011,
	14'b1100001100100,
	14'b1100001100101,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1110001010011,
	14'b1110001010100,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1111001010011,
	14'b1111001010100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b10000001010011,
	14'b10000001010100,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001010011,
	14'b10001001010100,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[186] <= 1'b1;
 		default: edge_mask_reg_p6[186] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100100,
	14'b1011001100101,
	14'b1011001100110,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1100001100100,
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1110001010100,
	14'b1110001010101,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1111001010100,
	14'b1111001010101,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001010100,
	14'b10000001010101,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10001001010100,
	14'b10001001010101,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[187] <= 1'b1;
 		default: edge_mask_reg_p6[187] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100101,
	14'b1011001100110,
	14'b1011001100111,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1110001010101,
	14'b1110001010110,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001010101,
	14'b1111001010110,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000001010101,
	14'b10000001010110,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001010101,
	14'b10001001010110,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000: edge_mask_reg_p6[188] <= 1'b1;
 		default: edge_mask_reg_p6[188] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100110,
	14'b1011001100111,
	14'b1011001101000,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101011110000,
	14'b1110001010110,
	14'b1110001010111,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1111001010110,
	14'b1111001010111,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010110,
	14'b10000001010111,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001001010110,
	14'b10001001010111,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010001110100,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[189] <= 1'b1;
 		default: edge_mask_reg_p6[189] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001100111,
	14'b1011001101000,
	14'b1011001101001,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001010111,
	14'b1110001011000,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100000,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110000,
	14'b1110010110110,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111001010111,
	14'b1111001011000,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010111,
	14'b10000001011000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10001001010111,
	14'b10001001011000,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[190] <= 1'b1;
 		default: edge_mask_reg_p6[190] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001101000,
	14'b1011001101001,
	14'b1011001101010,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011001111010,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001101010,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001101010,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110001011000,
	14'b1110001011001,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001101010,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110001111011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010001011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1111001011000,
	14'b1111001011001,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001101010,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111001111011,
	14'b1111010000001,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001011000,
	14'b10000001011001,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001101010,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000001111011,
	14'b10000010000001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001001011000,
	14'b10001001011001,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001101010,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001001111011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010001: edge_mask_reg_p6[191] <= 1'b1;
 		default: edge_mask_reg_p6[191] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110000,
	14'b1010010000000,
	14'b1010010010000,
	14'b1011001110000,
	14'b1011010000000,
	14'b1011010010000,
	14'b1100001110000,
	14'b1100010000000,
	14'b1100010010000,
	14'b1101001110000,
	14'b1101010000000,
	14'b1101010010000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010010100000,
	14'b10010010110000: edge_mask_reg_p6[192] <= 1'b1;
 		default: edge_mask_reg_p6[192] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110000,
	14'b1010001110001,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010010000,
	14'b1010010010001,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1110001100000,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010011000000: edge_mask_reg_p6[193] <= 1'b1;
 		default: edge_mask_reg_p6[193] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110000,
	14'b1010001110001,
	14'b1010001110010,
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1011001110000,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100001,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011010110000,
	14'b10011011000000: edge_mask_reg_p6[194] <= 1'b1;
 		default: edge_mask_reg_p6[194] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110001,
	14'b1010001110010,
	14'b1010001110011,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1011001110001,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100010,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10010010000000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011100000,
	14'b10100011100000,
	14'b10100011110000: edge_mask_reg_p6[195] <= 1'b1;
 		default: edge_mask_reg_p6[195] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010001110010,
	14'b1010001110011,
	14'b1010001110100,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1011001110010,
	14'b1011001110011,
	14'b1011001110100,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100011,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000001,
	14'b1111011000010,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[196] <= 1'b1;
 		default: edge_mask_reg_p6[196] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001110011,
	14'b1011001110100,
	14'b1011001110101,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100100,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000010,
	14'b1111011000011,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011110000,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[197] <= 1'b1;
 		default: edge_mask_reg_p6[197] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001110100,
	14'b1011001110101,
	14'b1011001110110,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100101,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011110000,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[198] <= 1'b1;
 		default: edge_mask_reg_p6[198] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001110101,
	14'b1011001110110,
	14'b1011001110111,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100110,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[199] <= 1'b1;
 		default: edge_mask_reg_p6[199] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001110110,
	14'b1011001110111,
	14'b1011001111000,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010000,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[200] <= 1'b1;
 		default: edge_mask_reg_p6[200] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001110111,
	14'b1011001111000,
	14'b1011001111001,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010101000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000: edge_mask_reg_p6[201] <= 1'b1;
 		default: edge_mask_reg_p6[201] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011001111000,
	14'b1011001111001,
	14'b1011001111010,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100011110000,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010001011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000110,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100001: edge_mask_reg_p6[202] <= 1'b1;
 		default: edge_mask_reg_p6[202] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000000,
	14'b1010010010000,
	14'b1010010100000,
	14'b1011010000000,
	14'b1011010010000,
	14'b1011010100000,
	14'b1100010000000,
	14'b1100010010000,
	14'b1100010100000,
	14'b1101010000000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010110000: edge_mask_reg_p6[203] <= 1'b1;
 		default: edge_mask_reg_p6[203] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010100000,
	14'b1010010100001,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10010010110000,
	14'b10010011000000: edge_mask_reg_p6[204] <= 1'b1;
 		default: edge_mask_reg_p6[204] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000000,
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1011010000000,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011011000000,
	14'b10011011010000: edge_mask_reg_p6[205] <= 1'b1;
 		default: edge_mask_reg_p6[205] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000001,
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1011010000001,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110010,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011010000: edge_mask_reg_p6[206] <= 1'b1;
 		default: edge_mask_reg_p6[206] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000010,
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1011010000010,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110011,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[207] <= 1'b1;
 		default: edge_mask_reg_p6[207] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010000011,
	14'b1010010000100,
	14'b1010010000101,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1011010000011,
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110100,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[208] <= 1'b1;
 		default: edge_mask_reg_p6[208] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010000100,
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110101,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010010,
	14'b1111011010011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[209] <= 1'b1;
 		default: edge_mask_reg_p6[209] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010000101,
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110110,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[210] <= 1'b1;
 		default: edge_mask_reg_p6[210] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010000110,
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110111,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[211] <= 1'b1;
 		default: edge_mask_reg_p6[211] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010000111,
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010111000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010000,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10101011010000,
	14'b10101011100000: edge_mask_reg_p6[212] <= 1'b1;
 		default: edge_mask_reg_p6[212] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010001000,
	14'b1011010001001,
	14'b1011010001010,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111001,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010011011,
	14'b1110010100000,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[213] <= 1'b1;
 		default: edge_mask_reg_p6[213] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010000,
	14'b1010010100000,
	14'b1010010110000,
	14'b1011010010000,
	14'b1011010100000,
	14'b1011010110000,
	14'b1100010010000,
	14'b1100010100000,
	14'b1100010110000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000: edge_mask_reg_p6[214] <= 1'b1;
 		default: edge_mask_reg_p6[214] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010110000,
	14'b1010010110001,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10010011000000,
	14'b10010011010000: edge_mask_reg_p6[215] <= 1'b1;
 		default: edge_mask_reg_p6[215] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010000,
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1011010010000,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000: edge_mask_reg_p6[216] <= 1'b1;
 		default: edge_mask_reg_p6[216] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010001,
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1011010010001,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000010,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000: edge_mask_reg_p6[217] <= 1'b1;
 		default: edge_mask_reg_p6[217] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010010,
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1011010010010,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000011,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010010,
	14'b1110011010011,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000: edge_mask_reg_p6[218] <= 1'b1;
 		default: edge_mask_reg_p6[218] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010010011,
	14'b1010010010100,
	14'b1010010010101,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1011010010011,
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000100,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[219] <= 1'b1;
 		default: edge_mask_reg_p6[219] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010010100,
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000101,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010010011,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[220] <= 1'b1;
 		default: edge_mask_reg_p6[220] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010010101,
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000110,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[221] <= 1'b1;
 		default: edge_mask_reg_p6[221] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010010110,
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000111,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000: edge_mask_reg_p6[222] <= 1'b1;
 		default: edge_mask_reg_p6[222] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010010111,
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011001000,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110101,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[223] <= 1'b1;
 		default: edge_mask_reg_p6[223] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010011000,
	14'b1011010011001,
	14'b1011010011010,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010101011,
	14'b1110010110000,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010: edge_mask_reg_p6[224] <= 1'b1;
 		default: edge_mask_reg_p6[224] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100000,
	14'b1010010110000,
	14'b1010011000000,
	14'b1011010100000,
	14'b1011010110000,
	14'b1011011000000,
	14'b1100010100000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001: edge_mask_reg_p6[225] <= 1'b1;
 		default: edge_mask_reg_p6[225] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010011000000,
	14'b1010011000001,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010011010000,
	14'b10010011100000: edge_mask_reg_p6[226] <= 1'b1;
 		default: edge_mask_reg_p6[226] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100000,
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1011010100000,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001: edge_mask_reg_p6[227] <= 1'b1;
 		default: edge_mask_reg_p6[227] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100001,
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1011010100001,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010010,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100001,
	14'b1110011100010,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011011010000,
	14'b10011011100000: edge_mask_reg_p6[228] <= 1'b1;
 		default: edge_mask_reg_p6[228] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100010,
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1011010100010,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010011,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100010,
	14'b1110011100011,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001: edge_mask_reg_p6[229] <= 1'b1;
 		default: edge_mask_reg_p6[229] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010100011,
	14'b1010010100100,
	14'b1010010100101,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1011010100011,
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010100,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100011,
	14'b1110011100100,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[230] <= 1'b1;
 		default: edge_mask_reg_p6[230] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010100100,
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010101,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100100,
	14'b1110011100101,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[231] <= 1'b1;
 		default: edge_mask_reg_p6[231] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010100101,
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010110,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[232] <= 1'b1;
 		default: edge_mask_reg_p6[232] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010100110,
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010111,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[233] <= 1'b1;
 		default: edge_mask_reg_p6[233] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010100111,
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011011000,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000: edge_mask_reg_p6[234] <= 1'b1;
 		default: edge_mask_reg_p6[234] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010101000,
	14'b1011010101001,
	14'b1011010101010,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110010111011,
	14'b1110011000000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010: edge_mask_reg_p6[235] <= 1'b1;
 		default: edge_mask_reg_p6[235] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110000,
	14'b1010011000000,
	14'b1010011010000,
	14'b1011010110000,
	14'b1011011000000,
	14'b1011011010000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001: edge_mask_reg_p6[236] <= 1'b1;
 		default: edge_mask_reg_p6[236] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110000,
	14'b1010010110001,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011010000,
	14'b1010011010001,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010011100000,
	14'b10010011110000: edge_mask_reg_p6[237] <= 1'b1;
 		default: edge_mask_reg_p6[237] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110000,
	14'b1010010110001,
	14'b1010010110010,
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1011010110000,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000: edge_mask_reg_p6[238] <= 1'b1;
 		default: edge_mask_reg_p6[238] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110001,
	14'b1010010110010,
	14'b1010010110011,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1011010110001,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10011011100000,
	14'b10011011110000: edge_mask_reg_p6[239] <= 1'b1;
 		default: edge_mask_reg_p6[239] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110010,
	14'b1010010110011,
	14'b1010010110100,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1011010110010,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001: edge_mask_reg_p6[240] <= 1'b1;
 		default: edge_mask_reg_p6[240] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110011,
	14'b1010010110100,
	14'b1010010110101,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1011010110011,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001: edge_mask_reg_p6[241] <= 1'b1;
 		default: edge_mask_reg_p6[241] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010010110100,
	14'b1010010110101,
	14'b1010010110110,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1011010110100,
	14'b1011010110101,
	14'b1011010110110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110100,
	14'b1110011110101,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[242] <= 1'b1;
 		default: edge_mask_reg_p6[242] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010110101,
	14'b1011010110110,
	14'b1011010110111,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[243] <= 1'b1;
 		default: edge_mask_reg_p6[243] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010110110,
	14'b1011010110111,
	14'b1011010111000,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110110,
	14'b1110011110111,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010110000,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[244] <= 1'b1;
 		default: edge_mask_reg_p6[244] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010110111,
	14'b1011010111000,
	14'b1011010111001,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011101000,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[245] <= 1'b1;
 		default: edge_mask_reg_p6[245] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011010111000,
	14'b1011010111001,
	14'b1011010111010,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101001,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011001011,
	14'b1110011010000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[246] <= 1'b1;
 		default: edge_mask_reg_p6[246] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000000,
	14'b1010011010000,
	14'b1010011100000,
	14'b1011011000000,
	14'b1011011010000,
	14'b1011011100000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001: edge_mask_reg_p6[247] <= 1'b1;
 		default: edge_mask_reg_p6[247] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011100000,
	14'b1010011100001,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10010011110000: edge_mask_reg_p6[248] <= 1'b1;
 		default: edge_mask_reg_p6[248] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000000,
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1011011000000,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000: edge_mask_reg_p6[249] <= 1'b1;
 		default: edge_mask_reg_p6[249] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000001,
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1011011000001,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000001,
	14'b1110100000010,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011011110000: edge_mask_reg_p6[250] <= 1'b1;
 		default: edge_mask_reg_p6[250] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000010,
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1011011000010,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000010,
	14'b1110100000011,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[251] <= 1'b1;
 		default: edge_mask_reg_p6[251] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000011,
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1011011000011,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000011,
	14'b1110100000100,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001: edge_mask_reg_p6[252] <= 1'b1;
 		default: edge_mask_reg_p6[252] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011000100,
	14'b1010011000101,
	14'b1010011000110,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1011011000100,
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[253] <= 1'b1;
 		default: edge_mask_reg_p6[253] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011000101,
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10010011000000,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011110000: edge_mask_reg_p6[254] <= 1'b1;
 		default: edge_mask_reg_p6[254] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011000110,
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011110000: edge_mask_reg_p6[255] <= 1'b1;
 		default: edge_mask_reg_p6[255] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011000111,
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011111000,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010110000,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000: edge_mask_reg_p6[256] <= 1'b1;
 		default: edge_mask_reg_p6[256] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011001000,
	14'b1011011001001,
	14'b1011011001010,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111001,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011011011,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[257] <= 1'b1;
 		default: edge_mask_reg_p6[257] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011010000,
	14'b1011011100000,
	14'b1011011110000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000: edge_mask_reg_p6[258] <= 1'b1;
 		default: edge_mask_reg_p6[258] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011110000,
	14'b1010011110001,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001: edge_mask_reg_p6[259] <= 1'b1;
 		default: edge_mask_reg_p6[259] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010000,
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1011011010000,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010011010000,
	14'b10010011110000,
	14'b10010100000000: edge_mask_reg_p6[260] <= 1'b1;
 		default: edge_mask_reg_p6[260] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010001,
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1011011010001,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000: edge_mask_reg_p6[261] <= 1'b1;
 		default: edge_mask_reg_p6[261] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010010,
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1011011010010,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[262] <= 1'b1;
 		default: edge_mask_reg_p6[262] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010011,
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1011011010011,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001: edge_mask_reg_p6[263] <= 1'b1;
 		default: edge_mask_reg_p6[263] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010100,
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1011011010100,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[264] <= 1'b1;
 		default: edge_mask_reg_p6[264] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011010101,
	14'b1010011010110,
	14'b1010011010111,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1011011010101,
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[265] <= 1'b1;
 		default: edge_mask_reg_p6[265] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011010110,
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10001011000000,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[266] <= 1'b1;
 		default: edge_mask_reg_p6[266] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011010111,
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100000,
	14'b10000011000000,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100000010: edge_mask_reg_p6[267] <= 1'b1;
 		default: edge_mask_reg_p6[267] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011011000,
	14'b1011011011001,
	14'b1011011011010,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011010000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000000,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[268] <= 1'b1;
 		default: edge_mask_reg_p6[268] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011100000,
	14'b1011011110000,
	14'b1011100000000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100100000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100100000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000: edge_mask_reg_p6[269] <= 1'b1;
 		default: edge_mask_reg_p6[269] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010100000000,
	14'b1010100000001,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011100000000,
	14'b1011100000001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001: edge_mask_reg_p6[270] <= 1'b1;
 		default: edge_mask_reg_p6[270] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100000,
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100000010,
	14'b1011011100000,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100000010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000: edge_mask_reg_p6[271] <= 1'b1;
 		default: edge_mask_reg_p6[271] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100001,
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100000011,
	14'b1011011100001,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100000011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001: edge_mask_reg_p6[272] <= 1'b1;
 		default: edge_mask_reg_p6[272] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100010,
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1011011100010,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000: edge_mask_reg_p6[273] <= 1'b1;
 		default: edge_mask_reg_p6[273] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100011,
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1011011100011,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001: edge_mask_reg_p6[274] <= 1'b1;
 		default: edge_mask_reg_p6[274] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100100,
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1011011100100,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[275] <= 1'b1;
 		default: edge_mask_reg_p6[275] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011100101,
	14'b1010011100110,
	14'b1010011100111,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100000111,
	14'b1011011100101,
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[276] <= 1'b1;
 		default: edge_mask_reg_p6[276] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011100110,
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b10000011010000,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10001011010000,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[277] <= 1'b1;
 		default: edge_mask_reg_p6[277] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011100111,
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1111011010000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100000,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101011110010,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100000010,
	14'b10101100010000: edge_mask_reg_p6[278] <= 1'b1;
 		default: edge_mask_reg_p6[278] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011101000,
	14'b1011011101001,
	14'b1011011101010,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1110011010000,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011100000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011101011,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100001011,
	14'b1110100010000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[279] <= 1'b1;
 		default: edge_mask_reg_p6[279] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100000000,
	14'b1011100010000,
	14'b1011100100000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100110000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100110000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100100000: edge_mask_reg_p6[280] <= 1'b1;
 		default: edge_mask_reg_p6[280] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110000,
	14'b1010011110001,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100010000,
	14'b1010100010001,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100010000,
	14'b1011100010001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001: edge_mask_reg_p6[281] <= 1'b1;
 		default: edge_mask_reg_p6[281] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110000,
	14'b1010011110001,
	14'b1010011110010,
	14'b1010100000000,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100010010,
	14'b1011011110000,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011100000000,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100010010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[282] <= 1'b1;
 		default: edge_mask_reg_p6[282] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110001,
	14'b1010011110010,
	14'b1010011110011,
	14'b1010100000001,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100010011,
	14'b1011011110001,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011100000001,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100010011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001: edge_mask_reg_p6[283] <= 1'b1;
 		default: edge_mask_reg_p6[283] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110010,
	14'b1010011110011,
	14'b1010011110100,
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100010100,
	14'b1011011110010,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100010100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[284] <= 1'b1;
 		default: edge_mask_reg_p6[284] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110011,
	14'b1010011110100,
	14'b1010011110101,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100010101,
	14'b1011011110011,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100010101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001: edge_mask_reg_p6[285] <= 1'b1;
 		default: edge_mask_reg_p6[285] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110100,
	14'b1010011110101,
	14'b1010011110110,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100010110,
	14'b1011011110100,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100010110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10010011100000,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[286] <= 1'b1;
 		default: edge_mask_reg_p6[286] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010011110101,
	14'b1010011110110,
	14'b1010011110111,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100000111,
	14'b1010100010101,
	14'b1010100010110,
	14'b1010100010111,
	14'b1011011110101,
	14'b1011011110110,
	14'b1011011110111,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100010111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110100000000: edge_mask_reg_p6[287] <= 1'b1;
 		default: edge_mask_reg_p6[287] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011110110,
	14'b1011011110111,
	14'b1011011111000,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100011000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000: edge_mask_reg_p6[288] <= 1'b1;
 		default: edge_mask_reg_p6[288] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011110111,
	14'b1011011111000,
	14'b1011011111001,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100011001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100000010,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[289] <= 1'b1;
 		default: edge_mask_reg_p6[289] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011011111000,
	14'b1011011111001,
	14'b1011011111010,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110011111011,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100001011,
	14'b1110100010000,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[290] <= 1'b1;
 		default: edge_mask_reg_p6[290] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100010000,
	14'b1010100100000,
	14'b1010100110000,
	14'b1011100010000,
	14'b1011100100000,
	14'b1011100110000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1101100110000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000: edge_mask_reg_p6[291] <= 1'b1;
 		default: edge_mask_reg_p6[291] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100110000,
	14'b1010100110001,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10010100000000: edge_mask_reg_p6[292] <= 1'b1;
 		default: edge_mask_reg_p6[292] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100010000,
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1011100010000,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[293] <= 1'b1;
 		default: edge_mask_reg_p6[293] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100010001,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1011100010001,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000001,
	14'b10001101000010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[294] <= 1'b1;
 		default: edge_mask_reg_p6[294] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100000010,
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100010010,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100100100,
	14'b1011100000010,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100010010,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011100110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000010,
	14'b10001101000011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[295] <= 1'b1;
 		default: edge_mask_reg_p6[295] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100000011,
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100010011,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100100101,
	14'b1011100000011,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100010011,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011100110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000011,
	14'b10001101000100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001: edge_mask_reg_p6[296] <= 1'b1;
 		default: edge_mask_reg_p6[296] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100000100,
	14'b1010100000101,
	14'b1010100000110,
	14'b1010100010100,
	14'b1010100010101,
	14'b1010100010110,
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100100110,
	14'b1011100000100,
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100010100,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100100110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[297] <= 1'b1;
 		default: edge_mask_reg_p6[297] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100000101,
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100010101,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100100111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110100000000: edge_mask_reg_p6[298] <= 1'b1;
 		default: edge_mask_reg_p6[298] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100000110,
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100010110,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100101000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000: edge_mask_reg_p6[299] <= 1'b1;
 		default: edge_mask_reg_p6[299] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100000111,
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100010111,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100101001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[300] <= 1'b1;
 		default: edge_mask_reg_p6[300] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100001000,
	14'b1011100001001,
	14'b1011100001010,
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100101010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[301] <= 1'b1;
 		default: edge_mask_reg_p6[301] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100000,
	14'b1010100110000,
	14'b1010101000000,
	14'b1011100100000,
	14'b1011100110000,
	14'b1011101000000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1101100100000,
	14'b1101100110000,
	14'b1101101000000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000: edge_mask_reg_p6[302] <= 1'b1;
 		default: edge_mask_reg_p6[302] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010101000000,
	14'b1010101000001,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1101100010000,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10010100000000,
	14'b10010100010000: edge_mask_reg_p6[303] <= 1'b1;
 		default: edge_mask_reg_p6[303] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100000,
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1011100100000,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[304] <= 1'b1;
 		default: edge_mask_reg_p6[304] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100001,
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1011100100001,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010001,
	14'b1111101010010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010001,
	14'b10000101010010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010001,
	14'b10001101010010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011100000000,
	14'b10011100010000: edge_mask_reg_p6[305] <= 1'b1;
 		default: edge_mask_reg_p6[305] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100010,
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1011100100010,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010010,
	14'b10001101010011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[306] <= 1'b1;
 		default: edge_mask_reg_p6[306] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100011,
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1011100100011,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010011,
	14'b10001101010100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001: edge_mask_reg_p6[307] <= 1'b1;
 		default: edge_mask_reg_p6[307] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100100100,
	14'b1010100100101,
	14'b1010100100110,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010100110110,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101000110,
	14'b1011100100100,
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010100,
	14'b10001101010101,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[308] <= 1'b1;
 		default: edge_mask_reg_p6[308] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100100101,
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110010,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[309] <= 1'b1;
 		default: edge_mask_reg_p6[309] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100100110,
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010110,
	14'b10001101010111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000100,
	14'b10010101000101,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[310] <= 1'b1;
 		default: edge_mask_reg_p6[310] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100100111,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000101,
	14'b10010101000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[311] <= 1'b1;
 		default: edge_mask_reg_p6[311] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100011000,
	14'b1011100011001,
	14'b1011100011010,
	14'b1011100101000,
	14'b1011100101001,
	14'b1011100101010,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011100111010,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100011011,
	14'b1110100100000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110000,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000001,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[312] <= 1'b1;
 		default: edge_mask_reg_p6[312] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110000,
	14'b1010101000000,
	14'b1010101010000,
	14'b1011100110000,
	14'b1011101000000,
	14'b1011101010000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1100101010000,
	14'b1101100110000,
	14'b1101101000000,
	14'b1101101010000,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000: edge_mask_reg_p6[313] <= 1'b1;
 		default: edge_mask_reg_p6[313] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110000,
	14'b1010100110001,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101010000,
	14'b1010101010001,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1101100100000,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[314] <= 1'b1;
 		default: edge_mask_reg_p6[314] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110000,
	14'b1010100110001,
	14'b1010100110010,
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1011100110000,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010101000000: edge_mask_reg_p6[315] <= 1'b1;
 		default: edge_mask_reg_p6[315] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110001,
	14'b1010100110010,
	14'b1010100110011,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1011100110001,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1101100100010,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100001,
	14'b1111101100010,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100001,
	14'b10000101100010,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100001,
	14'b10001101100010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[316] <= 1'b1;
 		default: edge_mask_reg_p6[316] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110010,
	14'b1010100110011,
	14'b1010100110100,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1011100110010,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1101100100011,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100010,
	14'b1111101100011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100010,
	14'b10000101100011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100010,
	14'b10001101100011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000: edge_mask_reg_p6[317] <= 1'b1;
 		default: edge_mask_reg_p6[317] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010100110011,
	14'b1010100110100,
	14'b1010100110101,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1011100110011,
	14'b1011100110100,
	14'b1011100110101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100011,
	14'b1111101100100,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100011,
	14'b10000101100100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100011,
	14'b10001101100100,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[318] <= 1'b1;
 		default: edge_mask_reg_p6[318] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100110100,
	14'b1011100110101,
	14'b1011100110110,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010011,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[319] <= 1'b1;
 		default: edge_mask_reg_p6[319] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100110101,
	14'b1011100110110,
	14'b1011100110111,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100101,
	14'b10001101100110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010011,
	14'b10010101010100,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[320] <= 1'b1;
 		default: edge_mask_reg_p6[320] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100110110,
	14'b1011100110111,
	14'b1011100111000,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100110,
	14'b10001101100111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010100,
	14'b10010101010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[321] <= 1'b1;
 		default: edge_mask_reg_p6[321] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100110111,
	14'b1011100111000,
	14'b1011100111001,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000001,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100111,
	14'b10001101101000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010101,
	14'b10010101010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[322] <= 1'b1;
 		default: edge_mask_reg_p6[322] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011100111000,
	14'b1011100111001,
	14'b1011100111010,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101001010,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100101011,
	14'b1110100110000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101101000,
	14'b10001101101001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010: edge_mask_reg_p6[323] <= 1'b1;
 		default: edge_mask_reg_p6[323] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000000,
	14'b1010101010000,
	14'b1010101100000,
	14'b1011101000000,
	14'b1011101010000,
	14'b1011101100000,
	14'b1100101000000,
	14'b1100101010000,
	14'b1100101100000,
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101100000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100110000: edge_mask_reg_p6[324] <= 1'b1;
 		default: edge_mask_reg_p6[324] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101100000,
	14'b1010101100001,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[325] <= 1'b1;
 		default: edge_mask_reg_p6[325] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000000,
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1011101000000,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101010000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[326] <= 1'b1;
 		default: edge_mask_reg_p6[326] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000001,
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1011101000001,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1101100110010,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110001,
	14'b1111101110010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110001,
	14'b10000101110010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110001,
	14'b10001101110010,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[327] <= 1'b1;
 		default: edge_mask_reg_p6[327] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000010,
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1011101000010,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1101100110011,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110010,
	14'b1111101110011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110010,
	14'b10000101110011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110010,
	14'b10001101110011,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000: edge_mask_reg_p6[328] <= 1'b1;
 		default: edge_mask_reg_p6[328] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101000011,
	14'b1010101000100,
	14'b1010101000101,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101100101,
	14'b1011101000011,
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1101100110100,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1111100010010,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110011,
	14'b1111101110100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110011,
	14'b10000101110100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110011,
	14'b10001101110100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[329] <= 1'b1;
 		default: edge_mask_reg_p6[329] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101000100,
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1101100110101,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1111100010011,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110100,
	14'b1111101110101,
	14'b10000011110000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110100,
	14'b10000101110101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110100,
	14'b10001101110101,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[330] <= 1'b1;
 		default: edge_mask_reg_p6[330] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101000101,
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1101100110110,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1111011110000,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110101,
	14'b1111101110110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110101,
	14'b10000101110110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110101,
	14'b10001101110110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000: edge_mask_reg_p6[331] <= 1'b1;
 		default: edge_mask_reg_p6[331] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101000110,
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1110011110000,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010100,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110110,
	14'b10001101110111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[332] <= 1'b1;
 		default: edge_mask_reg_p6[332] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101000111,
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110111,
	14'b10001101111000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[333] <= 1'b1;
 		default: edge_mask_reg_p6[333] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101001000,
	14'b1011101001001,
	14'b1011101001010,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110100111011,
	14'b1110101000000,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101111000,
	14'b10001101111001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010101,
	14'b10010101010110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[334] <= 1'b1;
 		default: edge_mask_reg_p6[334] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010000,
	14'b1010101100000,
	14'b1010101110000,
	14'b1011101010000,
	14'b1011101100000,
	14'b1011101110000,
	14'b1100101010000,
	14'b1100101100000,
	14'b1100101110000,
	14'b1101101010000,
	14'b1101101100000,
	14'b1101101110000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10010100110000,
	14'b10010101000000: edge_mask_reg_p6[335] <= 1'b1;
 		default: edge_mask_reg_p6[335] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101110000,
	14'b1010101110001,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001: edge_mask_reg_p6[336] <= 1'b1;
 		default: edge_mask_reg_p6[336] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010000,
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1011101010000,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[337] <= 1'b1;
 		default: edge_mask_reg_p6[337] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010001,
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1011101010001,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1101101000010,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000001,
	14'b1111110000010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000001,
	14'b10000110000010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000001,
	14'b10001110000010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000: edge_mask_reg_p6[338] <= 1'b1;
 		default: edge_mask_reg_p6[338] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010010,
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010101110100,
	14'b1011101010010,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1101101000011,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000010,
	14'b1111110000011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000010,
	14'b10000110000011,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000010,
	14'b10001110000011,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[339] <= 1'b1;
 		default: edge_mask_reg_p6[339] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101010011,
	14'b1010101010100,
	14'b1010101010101,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101100101,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010101110101,
	14'b1011101010011,
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1101101000100,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000011,
	14'b1111110000100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000011,
	14'b10000110000100,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000011,
	14'b10001110000100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100001,
	14'b10010101100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[340] <= 1'b1;
 		default: edge_mask_reg_p6[340] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101010100,
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1101101000101,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000100,
	14'b1111110000101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000100,
	14'b10000110000101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000100,
	14'b10001110000101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[341] <= 1'b1;
 		default: edge_mask_reg_p6[341] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101010101,
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1101101000110,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000101,
	14'b1111110000110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000101,
	14'b10000110000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000101,
	14'b10001110000110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[342] <= 1'b1;
 		default: edge_mask_reg_p6[342] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101010110,
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1101101000111,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000110,
	14'b1111110000111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000110,
	14'b10000110000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010000,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000110,
	14'b10001110000111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101010000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[343] <= 1'b1;
 		default: edge_mask_reg_p6[343] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101010111,
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000111,
	14'b1111110001000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000111,
	14'b10000110001000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000111,
	14'b10001110001000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10101100100000: edge_mask_reg_p6[344] <= 1'b1;
 		default: edge_mask_reg_p6[344] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101011000,
	14'b1011101011001,
	14'b1011101011010,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100110000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101000000,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101001011,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110001000,
	14'b1110110001001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110001000,
	14'b10001110001001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010100,
	14'b10010101010101,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[345] <= 1'b1;
 		default: edge_mask_reg_p6[345] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100000,
	14'b1010101110000,
	14'b1010110000000,
	14'b1011101100000,
	14'b1011101110000,
	14'b1011110000000,
	14'b1100101100000,
	14'b1100101110000,
	14'b1100110000000,
	14'b1101101100000,
	14'b1101101110000,
	14'b1101110000000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10010101000000,
	14'b10010101010000: edge_mask_reg_p6[346] <= 1'b1;
 		default: edge_mask_reg_p6[346] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010110000000,
	14'b1010110000001,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011110000000,
	14'b1011110000001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110000001,
	14'b1101101010000,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110010000,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110010000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001: edge_mask_reg_p6[347] <= 1'b1;
 		default: edge_mask_reg_p6[347] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100000,
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110000010,
	14'b1011101100000,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110000010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100110000,
	14'b10011101000000: edge_mask_reg_p6[348] <= 1'b1;
 		default: edge_mask_reg_p6[348] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100001,
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110000011,
	14'b1011101100001,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110000011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1101101010010,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010001,
	14'b1110110010010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010001,
	14'b10000110010010,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[349] <= 1'b1;
 		default: edge_mask_reg_p6[349] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101100010,
	14'b1010101100011,
	14'b1010101100100,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010101110100,
	14'b1010110000010,
	14'b1010110000011,
	14'b1010110000100,
	14'b1011101100010,
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110000100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1101101010011,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010010,
	14'b1110110010011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010010,
	14'b1111110010011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010010,
	14'b10000110010011,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010010,
	14'b10001110010011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[350] <= 1'b1;
 		default: edge_mask_reg_p6[350] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101100011,
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110000101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1101101010100,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010011,
	14'b1110110010100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010011,
	14'b1111110010100,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010011,
	14'b10000110010100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010011,
	14'b10001110010100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110001,
	14'b10010101110010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[351] <= 1'b1;
 		default: edge_mask_reg_p6[351] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101100100,
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110000110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1101101010101,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010100,
	14'b1110110010101,
	14'b1111100000000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010100,
	14'b1111110010101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010100,
	14'b10000110010101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010100,
	14'b10001110010101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110010,
	14'b10010101110011,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[352] <= 1'b1;
 		default: edge_mask_reg_p6[352] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101100101,
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110000111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1101101010110,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1110100000000,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010101,
	14'b1110110010110,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010101,
	14'b1111110010110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010101,
	14'b10000110010110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010101,
	14'b10001110010110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001,
	14'b10101101000000: edge_mask_reg_p6[353] <= 1'b1;
 		default: edge_mask_reg_p6[353] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101100110,
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110001000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1101101010111,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010110,
	14'b1110110010111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010110,
	14'b1111110010111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010110,
	14'b10000110010111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010110,
	14'b10001110010111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[354] <= 1'b1;
 		default: edge_mask_reg_p6[354] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101100111,
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110001001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101011000,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010111,
	14'b1110110011000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010111,
	14'b1111110011000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010111,
	14'b10000110011000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010111,
	14'b10001110011000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010: edge_mask_reg_p6[355] <= 1'b1;
 		default: edge_mask_reg_p6[355] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101101000,
	14'b1011101101001,
	14'b1011101101010,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110001010,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101101011001,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101011011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110101111011,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110011000,
	14'b1110110011001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110011000,
	14'b1111110011001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110011000,
	14'b10000110011001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110011000,
	14'b10001110011001,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010: edge_mask_reg_p6[356] <= 1'b1;
 		default: edge_mask_reg_p6[356] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110000,
	14'b1010110000000,
	14'b1010110010000,
	14'b1011101110000,
	14'b1011110000000,
	14'b1011110010000,
	14'b1100101110000,
	14'b1100110000000,
	14'b1100110010000,
	14'b1101101110000,
	14'b1101110000000,
	14'b1101110010000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110010000,
	14'b1111101010000,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000101010000,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001101010000,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110010000,
	14'b10010101010000,
	14'b10010101100000: edge_mask_reg_p6[357] <= 1'b1;
 		default: edge_mask_reg_p6[357] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110000,
	14'b1010101110001,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110010000,
	14'b1010110010001,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110010000,
	14'b1011110010001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110010000,
	14'b1100110010001,
	14'b1101101100000,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110010000,
	14'b1101110010001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110100000,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10001110010001,
	14'b10010101000000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011101000000: edge_mask_reg_p6[358] <= 1'b1;
 		default: edge_mask_reg_p6[358] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110000,
	14'b1010101110001,
	14'b1010101110010,
	14'b1010110000000,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110010000,
	14'b1010110010001,
	14'b1010110010010,
	14'b1011101110000,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011110000000,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110010000,
	14'b1011110010001,
	14'b1011110010010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110010000,
	14'b1100110010001,
	14'b1100110010010,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110010000,
	14'b1101110010001,
	14'b1101110010010,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110100000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110100000,
	14'b1111110100001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10000110100001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110100000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10011100010000,
	14'b10011101000000,
	14'b10011101010000,
	14'b10100100010000: edge_mask_reg_p6[359] <= 1'b1;
 		default: edge_mask_reg_p6[359] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1010101110001,
	14'b1010101110010,
	14'b1010101110011,
	14'b1010110000001,
	14'b1010110000010,
	14'b1010110000011,
	14'b1010110010001,
	14'b1010110010010,
	14'b1010110010011,
	14'b1011101110001,
	14'b1011101110010,
	14'b1011101110011,
	14'b1011110000001,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110010001,
	14'b1011110010010,
	14'b1011110010011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110010001,
	14'b1100110010010,
	14'b1100110010011,
	14'b1101101100010,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110010011,
	14'b1110101010010,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110100001,
	14'b1110110100010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110100001,
	14'b1111110100010,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110100001,
	14'b10000110100010,
	14'b10001100010000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110100001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101100010000: edge_mask_reg_p6[360] <= 1'b1;
 		default: edge_mask_reg_p6[360] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110010,
	14'b1011101110011,
	14'b1011101110100,
	14'b1011110000010,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110010010,
	14'b1011110010011,
	14'b1011110010100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110010010,
	14'b1100110010011,
	14'b1100110010100,
	14'b1101101100011,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110010100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110100010,
	14'b1110110100011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110100010,
	14'b1111110100011,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110100010,
	14'b10000110100011,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110100010,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[361] <= 1'b1;
 		default: edge_mask_reg_p6[361] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110011,
	14'b1011101110100,
	14'b1011101110101,
	14'b1011110000011,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110010011,
	14'b1011110010100,
	14'b1011110010101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110010011,
	14'b1100110010100,
	14'b1100110010101,
	14'b1101101100100,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110010101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110100011,
	14'b1110110100100,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110100011,
	14'b1111110100100,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110100011,
	14'b10000110100100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110100011,
	14'b10001110100100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000001,
	14'b10010110000010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[362] <= 1'b1;
 		default: edge_mask_reg_p6[362] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110100,
	14'b1011101110101,
	14'b1011101110110,
	14'b1011110000100,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110010100,
	14'b1011110010101,
	14'b1011110010110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110010100,
	14'b1100110010101,
	14'b1100110010110,
	14'b1101101100101,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110010110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110100100,
	14'b1110110100101,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110100100,
	14'b1111110100101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110100100,
	14'b10000110100101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110100100,
	14'b10001110100101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000010,
	14'b10010110000011,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[363] <= 1'b1;
 		default: edge_mask_reg_p6[363] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110101,
	14'b1011101110110,
	14'b1011101110111,
	14'b1011110000101,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110010101,
	14'b1011110010110,
	14'b1011110010111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110010101,
	14'b1100110010110,
	14'b1100110010111,
	14'b1101101100110,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110010111,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110100101,
	14'b1110110100110,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110100101,
	14'b1111110100110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110100101,
	14'b10000110100110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110100101,
	14'b10001110100110,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000011,
	14'b10010110000100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[364] <= 1'b1;
 		default: edge_mask_reg_p6[364] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110110,
	14'b1011101110111,
	14'b1011101111000,
	14'b1011110000110,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110010110,
	14'b1011110010111,
	14'b1011110011000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110010110,
	14'b1100110010111,
	14'b1100110011000,
	14'b1101100000000,
	14'b1101101100111,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110011000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110100110,
	14'b1110110100111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110100110,
	14'b1111110100111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110100110,
	14'b10000110100111,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110100110,
	14'b10001110100111,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[365] <= 1'b1;
 		default: edge_mask_reg_p6[365] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101110111,
	14'b1011101111000,
	14'b1011101111001,
	14'b1011110000111,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110010111,
	14'b1011110011000,
	14'b1011110011001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110010111,
	14'b1100110011000,
	14'b1100110011001,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101101000,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110011001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100001,
	14'b1110101000000,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010000,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110100111,
	14'b1110110101000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110100111,
	14'b1111110101000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110100111,
	14'b10000110101000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110100111,
	14'b10001110101000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[366] <= 1'b1;
 		default: edge_mask_reg_p6[366] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1011101111000,
	14'b1011101111001,
	14'b1011101111010,
	14'b1011110001000,
	14'b1011110001001,
	14'b1011110001010,
	14'b1011110011000,
	14'b1011110011001,
	14'b1011110011010,
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1100110011000,
	14'b1100110011001,
	14'b1100110011010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101101001,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110011000,
	14'b1101110011001,
	14'b1101110011010,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101101011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110101111011,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110001011,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110011010,
	14'b1110110101000,
	14'b1110110101001,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110000,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110001011,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110011010,
	14'b1111110101000,
	14'b1111110101001,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110000,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110001011,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110011010,
	14'b10000110101000,
	14'b10000110101001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110001011,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110011010,
	14'b10001110101000,
	14'b10001110101001,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010: edge_mask_reg_p6[367] <= 1'b1;
 		default: edge_mask_reg_p6[367] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100000,
	14'b1100001110000,
	14'b1100010000000,
	14'b1101001100000,
	14'b1101001110000,
	14'b1101010000000,
	14'b1110001100000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10010001100000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10011010010000,
	14'b10011010100000: edge_mask_reg_p6[368] <= 1'b1;
 		default: edge_mask_reg_p6[368] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100000,
	14'b1100001100001,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1111001010000,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b10000001010000,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001010000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010110000: edge_mask_reg_p6[369] <= 1'b1;
 		default: edge_mask_reg_p6[369] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100000,
	14'b1100001100001,
	14'b1100001100010,
	14'b1100001110000,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1111001010000,
	14'b1111001010001,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b10000001010000,
	14'b10000001010001,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10001001010000,
	14'b10001001010001,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10010001010000,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001: edge_mask_reg_p6[370] <= 1'b1;
 		default: edge_mask_reg_p6[370] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100001,
	14'b1100001100010,
	14'b1100001100011,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1111001010001,
	14'b1111001010010,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100001,
	14'b1111010100010,
	14'b10000001010001,
	14'b10000001010010,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10001001010001,
	14'b10001001010010,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001010001,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011001110000,
	14'b10011010000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100011100000,
	14'b10100011110000: edge_mask_reg_p6[371] <= 1'b1;
 		default: edge_mask_reg_p6[371] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100010,
	14'b1100001100011,
	14'b1100001100100,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1111001010010,
	14'b1111001010011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100010,
	14'b1111010100011,
	14'b10000001010010,
	14'b10000001010011,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10001001010010,
	14'b10001001010011,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011100000,
	14'b10010001010010,
	14'b10010001010011,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10101011100000: edge_mask_reg_p6[372] <= 1'b1;
 		default: edge_mask_reg_p6[372] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100011,
	14'b1100001100100,
	14'b1100001100101,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1111001010011,
	14'b1111001010100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b10000001010011,
	14'b10000001010100,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001010011,
	14'b10001001010100,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010001010011,
	14'b10010001010100,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[373] <= 1'b1;
 		default: edge_mask_reg_p6[373] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100100,
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1111001010100,
	14'b1111001010101,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001010100,
	14'b10000001010101,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001010100,
	14'b10001001010101,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010001010100,
	14'b10010001010101,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011001110010,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[374] <= 1'b1;
 		default: edge_mask_reg_p6[374] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100101,
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110011110000,
	14'b1111001010101,
	14'b1111001010110,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110100,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001010101,
	14'b10000001010110,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001010101,
	14'b10001001010110,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010001010101,
	14'b10010001010110,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[375] <= 1'b1;
 		default: edge_mask_reg_p6[375] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100110,
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001010110,
	14'b1111001010111,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010110,
	14'b10000001010111,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001010110,
	14'b10001001010111,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001010110,
	14'b10010001010111,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010010000,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101011010000: edge_mask_reg_p6[376] <= 1'b1;
 		default: edge_mask_reg_p6[376] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001100111,
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111001010111,
	14'b1111001011000,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010111,
	14'b10000001011000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10001001010111,
	14'b10001001011000,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10010001010111,
	14'b10010001011000,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[377] <= 1'b1;
 		default: edge_mask_reg_p6[377] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001101000,
	14'b1100001101001,
	14'b1100001101010,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001101010,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001101010,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1111001011000,
	14'b1111001011001,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001101010,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111001111011,
	14'b1111010000001,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001011000,
	14'b10000001011001,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001101010,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000001111011,
	14'b10000010000001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001001011000,
	14'b10001001011001,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001101010,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001001111011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010001011000,
	14'b10010001011001,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001101010,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010001111011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010001011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001: edge_mask_reg_p6[378] <= 1'b1;
 		default: edge_mask_reg_p6[378] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110000,
	14'b1100010000000,
	14'b1100010010000,
	14'b1101001110000,
	14'b1101010000000,
	14'b1101010010000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010010000,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010001110000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000: edge_mask_reg_p6[379] <= 1'b1;
 		default: edge_mask_reg_p6[379] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110000,
	14'b1100001110001,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011011000000: edge_mask_reg_p6[380] <= 1'b1;
 		default: edge_mask_reg_p6[380] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110000,
	14'b1100001110001,
	14'b1100001110010,
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001100000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000: edge_mask_reg_p6[381] <= 1'b1;
 		default: edge_mask_reg_p6[381] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110001,
	14'b1100001110010,
	14'b1100001110011,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110001,
	14'b1111010110010,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010001100001,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011010000000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001: edge_mask_reg_p6[382] <= 1'b1;
 		default: edge_mask_reg_p6[382] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110010,
	14'b1100001110011,
	14'b1100001110100,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[383] <= 1'b1;
 		default: edge_mask_reg_p6[383] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110011,
	14'b1100001110100,
	14'b1100001110101,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[384] <= 1'b1;
 		default: edge_mask_reg_p6[384] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110100,
	14'b1100001110101,
	14'b1100001110110,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[385] <= 1'b1;
 		default: edge_mask_reg_p6[385] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110101,
	14'b1100001110110,
	14'b1100001110111,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[386] <= 1'b1;
 		default: edge_mask_reg_p6[386] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110110,
	14'b1100001110111,
	14'b1100001111000,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010000,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010010000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[387] <= 1'b1;
 		default: edge_mask_reg_p6[387] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001110111,
	14'b1100001111000,
	14'b1100001111001,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101011110000,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000101,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000: edge_mask_reg_p6[388] <= 1'b1;
 		default: edge_mask_reg_p6[388] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100001111000,
	14'b1100001111001,
	14'b1100001111010,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100000,
	14'b1110010101001,
	14'b1110010110000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010001011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010001011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001: edge_mask_reg_p6[389] <= 1'b1;
 		default: edge_mask_reg_p6[389] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000000,
	14'b1100010010000,
	14'b1100010100000,
	14'b1101010000000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010000000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000: edge_mask_reg_p6[390] <= 1'b1;
 		default: edge_mask_reg_p6[390] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10011010110000,
	14'b10011011000000: edge_mask_reg_p6[391] <= 1'b1;
 		default: edge_mask_reg_p6[391] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000000,
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010001110000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000: edge_mask_reg_p6[392] <= 1'b1;
 		default: edge_mask_reg_p6[392] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000001,
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001: edge_mask_reg_p6[393] <= 1'b1;
 		default: edge_mask_reg_p6[393] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000010,
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10100011000000,
	14'b10100011010000: edge_mask_reg_p6[394] <= 1'b1;
 		default: edge_mask_reg_p6[394] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000011,
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110100,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011110000: edge_mask_reg_p6[395] <= 1'b1;
 		default: edge_mask_reg_p6[395] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000100,
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110101,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[396] <= 1'b1;
 		default: edge_mask_reg_p6[396] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000101,
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110110,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011110000,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[397] <= 1'b1;
 		default: edge_mask_reg_p6[397] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000110,
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110111,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[398] <= 1'b1;
 		default: edge_mask_reg_p6[398] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010000111,
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010111000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011010000,
	14'b10101011100000: edge_mask_reg_p6[399] <= 1'b1;
 		default: edge_mask_reg_p6[399] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010001000,
	14'b1100010001001,
	14'b1100010001010,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110000,
	14'b1110010111001,
	14'b1110011000000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010011011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[400] <= 1'b1;
 		default: edge_mask_reg_p6[400] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010000,
	14'b1100010100000,
	14'b1100010110000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001: edge_mask_reg_p6[401] <= 1'b1;
 		default: edge_mask_reg_p6[401] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10011011000000,
	14'b10011011010000: edge_mask_reg_p6[402] <= 1'b1;
 		default: edge_mask_reg_p6[402] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010000,
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000: edge_mask_reg_p6[403] <= 1'b1;
 		default: edge_mask_reg_p6[403] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010001,
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000010,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000: edge_mask_reg_p6[404] <= 1'b1;
 		default: edge_mask_reg_p6[404] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010010,
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000011,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10100011010000: edge_mask_reg_p6[405] <= 1'b1;
 		default: edge_mask_reg_p6[405] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010011,
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000100,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[406] <= 1'b1;
 		default: edge_mask_reg_p6[406] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010100,
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000101,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100010,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[407] <= 1'b1;
 		default: edge_mask_reg_p6[407] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010101,
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000110,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10110011100000: edge_mask_reg_p6[408] <= 1'b1;
 		default: edge_mask_reg_p6[408] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010110,
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000111,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100000,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[409] <= 1'b1;
 		default: edge_mask_reg_p6[409] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010010111,
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011001000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[410] <= 1'b1;
 		default: edge_mask_reg_p6[410] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010011000,
	14'b1100010011001,
	14'b1100010011010,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011000000,
	14'b1110011001001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010101011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011001011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010: edge_mask_reg_p6[411] <= 1'b1;
 		default: edge_mask_reg_p6[411] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100000,
	14'b1100010110000,
	14'b1100011000000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001: edge_mask_reg_p6[412] <= 1'b1;
 		default: edge_mask_reg_p6[412] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10011011010000,
	14'b10011011100000: edge_mask_reg_p6[413] <= 1'b1;
 		default: edge_mask_reg_p6[413] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100000,
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000: edge_mask_reg_p6[414] <= 1'b1;
 		default: edge_mask_reg_p6[414] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100001,
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010010,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001: edge_mask_reg_p6[415] <= 1'b1;
 		default: edge_mask_reg_p6[415] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100010,
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010011,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000: edge_mask_reg_p6[416] <= 1'b1;
 		default: edge_mask_reg_p6[416] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100011,
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010100,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000: edge_mask_reg_p6[417] <= 1'b1;
 		default: edge_mask_reg_p6[417] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100100,
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010101,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101100000000: edge_mask_reg_p6[418] <= 1'b1;
 		default: edge_mask_reg_p6[418] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100101,
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010110,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010100011,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000: edge_mask_reg_p6[419] <= 1'b1;
 		default: edge_mask_reg_p6[419] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100110,
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010111,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000100,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111100000000,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[420] <= 1'b1;
 		default: edge_mask_reg_p6[420] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010100111,
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011011000,
	14'b1110100000000,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[421] <= 1'b1;
 		default: edge_mask_reg_p6[421] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010101000,
	14'b1100010101001,
	14'b1100010101010,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011011001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111010111011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011001011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001: edge_mask_reg_p6[422] <= 1'b1;
 		default: edge_mask_reg_p6[422] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110000,
	14'b1100011000000,
	14'b1100011010000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001: edge_mask_reg_p6[423] <= 1'b1;
 		default: edge_mask_reg_p6[423] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110000,
	14'b1100010110001,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000: edge_mask_reg_p6[424] <= 1'b1;
 		default: edge_mask_reg_p6[424] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110000,
	14'b1100010110001,
	14'b1100010110010,
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10011011100000,
	14'b10011011110000: edge_mask_reg_p6[425] <= 1'b1;
 		default: edge_mask_reg_p6[425] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110001,
	14'b1100010110010,
	14'b1100010110011,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100010,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001: edge_mask_reg_p6[426] <= 1'b1;
 		default: edge_mask_reg_p6[426] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110010,
	14'b1100010110011,
	14'b1100010110100,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100011,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110010,
	14'b1111011110011,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010: edge_mask_reg_p6[427] <= 1'b1;
 		default: edge_mask_reg_p6[427] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110011,
	14'b1100010110100,
	14'b1100010110101,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100100,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110011,
	14'b1111011110100,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000: edge_mask_reg_p6[428] <= 1'b1;
 		default: edge_mask_reg_p6[428] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110100,
	14'b1100010110101,
	14'b1100010110110,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100101,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110100,
	14'b1111011110101,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[429] <= 1'b1;
 		default: edge_mask_reg_p6[429] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110101,
	14'b1100010110110,
	14'b1100010110111,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100110,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[430] <= 1'b1;
 		default: edge_mask_reg_p6[430] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110110,
	14'b1100010110111,
	14'b1100010111000,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100111,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011010110000,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[431] <= 1'b1;
 		default: edge_mask_reg_p6[431] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010110111,
	14'b1100010111000,
	14'b1100010111001,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011101000,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[432] <= 1'b1;
 		default: edge_mask_reg_p6[432] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100010111000,
	14'b1100010111001,
	14'b1100010111010,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011101001,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011001011,
	14'b1111011010000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011011011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[433] <= 1'b1;
 		default: edge_mask_reg_p6[433] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000000,
	14'b1100011010000,
	14'b1100011100000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001: edge_mask_reg_p6[434] <= 1'b1;
 		default: edge_mask_reg_p6[434] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000: edge_mask_reg_p6[435] <= 1'b1;
 		default: edge_mask_reg_p6[435] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000000,
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[436] <= 1'b1;
 		default: edge_mask_reg_p6[436] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000001,
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110010,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001: edge_mask_reg_p6[437] <= 1'b1;
 		default: edge_mask_reg_p6[437] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000010,
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000010,
	14'b1111100000011,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010: edge_mask_reg_p6[438] <= 1'b1;
 		default: edge_mask_reg_p6[438] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000011,
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000011,
	14'b1111100000100,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100011100000,
	14'b10100011110000: edge_mask_reg_p6[439] <= 1'b1;
 		default: edge_mask_reg_p6[439] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000100,
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000: edge_mask_reg_p6[440] <= 1'b1;
 		default: edge_mask_reg_p6[440] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000101,
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110110,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011110000: edge_mask_reg_p6[441] <= 1'b1;
 		default: edge_mask_reg_p6[441] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000110,
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110111,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010000,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[442] <= 1'b1;
 		default: edge_mask_reg_p6[442] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011000111,
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011111000,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010110000,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000: edge_mask_reg_p6[443] <= 1'b1;
 		default: edge_mask_reg_p6[443] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011001000,
	14'b1100011001001,
	14'b1100011001010,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011111001,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011011011,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011101011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[444] <= 1'b1;
 		default: edge_mask_reg_p6[444] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010000,
	14'b1100011100000,
	14'b1100011110000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000: edge_mask_reg_p6[445] <= 1'b1;
 		default: edge_mask_reg_p6[445] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001: edge_mask_reg_p6[446] <= 1'b1;
 		default: edge_mask_reg_p6[446] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010000,
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011100000000: edge_mask_reg_p6[447] <= 1'b1;
 		default: edge_mask_reg_p6[447] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010001,
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000: edge_mask_reg_p6[448] <= 1'b1;
 		default: edge_mask_reg_p6[448] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010010,
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001: edge_mask_reg_p6[449] <= 1'b1;
 		default: edge_mask_reg_p6[449] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010011,
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[450] <= 1'b1;
 		default: edge_mask_reg_p6[450] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010100,
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000: edge_mask_reg_p6[451] <= 1'b1;
 		default: edge_mask_reg_p6[451] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010101,
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100100000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[452] <= 1'b1;
 		default: edge_mask_reg_p6[452] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010110,
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000111,
	14'b1110100001000,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10001011000000,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[453] <= 1'b1;
 		default: edge_mask_reg_p6[453] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011010111,
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100001000,
	14'b1110100001001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010000,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b10000011000000,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[454] <= 1'b1;
 		default: edge_mask_reg_p6[454] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011011000,
	14'b1100011011001,
	14'b1100011011010,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100000000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1111011000000,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[455] <= 1'b1;
 		default: edge_mask_reg_p6[455] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100000,
	14'b1100011110000,
	14'b1100100000000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100100000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000: edge_mask_reg_p6[456] <= 1'b1;
 		default: edge_mask_reg_p6[456] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001: edge_mask_reg_p6[457] <= 1'b1;
 		default: edge_mask_reg_p6[457] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011100000,
	14'b10011100010000: edge_mask_reg_p6[458] <= 1'b1;
 		default: edge_mask_reg_p6[458] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100001,
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001: edge_mask_reg_p6[459] <= 1'b1;
 		default: edge_mask_reg_p6[459] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100010,
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010: edge_mask_reg_p6[460] <= 1'b1;
 		default: edge_mask_reg_p6[460] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100011,
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[461] <= 1'b1;
 		default: edge_mask_reg_p6[461] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100100,
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000: edge_mask_reg_p6[462] <= 1'b1;
 		default: edge_mask_reg_p6[462] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100101,
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[463] <= 1'b1;
 		default: edge_mask_reg_p6[463] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100110,
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10001011010000,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10010011010000,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[464] <= 1'b1;
 		default: edge_mask_reg_p6[464] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100111,
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100011000,
	14'b1110100011001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b10000011010000,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[465] <= 1'b1;
 		default: edge_mask_reg_p6[465] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011101000,
	14'b1100011101001,
	14'b1100011101010,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100010000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100100000,
	14'b1111011010000,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011101011,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100001011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[466] <= 1'b1;
 		default: edge_mask_reg_p6[466] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000000,
	14'b1100100010000,
	14'b1100100100000,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110100100000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100110000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000: edge_mask_reg_p6[467] <= 1'b1;
 		default: edge_mask_reg_p6[467] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100011110001,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001: edge_mask_reg_p6[468] <= 1'b1;
 		default: edge_mask_reg_p6[468] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100011110001,
	14'b1100011110010,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011110000: edge_mask_reg_p6[469] <= 1'b1;
 		default: edge_mask_reg_p6[469] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110001,
	14'b1100011110010,
	14'b1100011110011,
	14'b1100100000001,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[470] <= 1'b1;
 		default: edge_mask_reg_p6[470] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110010,
	14'b1100011110011,
	14'b1100011110100,
	14'b1100100000010,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010: edge_mask_reg_p6[471] <= 1'b1;
 		default: edge_mask_reg_p6[471] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110011,
	14'b1100011110100,
	14'b1100011110101,
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[472] <= 1'b1;
 		default: edge_mask_reg_p6[472] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110100,
	14'b1100011110101,
	14'b1100011110110,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10010011100000,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10011011100000,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001: edge_mask_reg_p6[473] <= 1'b1;
 		default: edge_mask_reg_p6[473] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110101,
	14'b1100011110110,
	14'b1100011110111,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110100000000: edge_mask_reg_p6[474] <= 1'b1;
 		default: edge_mask_reg_p6[474] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110110,
	14'b1100011110111,
	14'b1100011111000,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[475] <= 1'b1;
 		default: edge_mask_reg_p6[475] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110111,
	14'b1100011111000,
	14'b1100011111001,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[476] <= 1'b1;
 		default: edge_mask_reg_p6[476] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011111000,
	14'b1100011111001,
	14'b1100011111010,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111011111011,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100001011,
	14'b1111100010000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100001011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[477] <= 1'b1;
 		default: edge_mask_reg_p6[477] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100010000,
	14'b1100100100000,
	14'b1100100110000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1101100110000,
	14'b1110100010000,
	14'b1110100100000,
	14'b1110100110000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000: edge_mask_reg_p6[478] <= 1'b1;
 		default: edge_mask_reg_p6[478] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000: edge_mask_reg_p6[479] <= 1'b1;
 		default: edge_mask_reg_p6[479] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100010000,
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011110000,
	14'b10011100000000: edge_mask_reg_p6[480] <= 1'b1;
 		default: edge_mask_reg_p6[480] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100010001,
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[481] <= 1'b1;
 		default: edge_mask_reg_p6[481] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100010010,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000010,
	14'b10010101000011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001: edge_mask_reg_p6[482] <= 1'b1;
 		default: edge_mask_reg_p6[482] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000011,
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100010011,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110001,
	14'b10011100110010,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[483] <= 1'b1;
 		default: edge_mask_reg_p6[483] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000100,
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100010100,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000: edge_mask_reg_p6[484] <= 1'b1;
 		default: edge_mask_reg_p6[484] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000101,
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100010101,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110100000000: edge_mask_reg_p6[485] <= 1'b1;
 		default: edge_mask_reg_p6[485] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000110,
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100010110,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[486] <= 1'b1;
 		default: edge_mask_reg_p6[486] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100000111,
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100010111,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[487] <= 1'b1;
 		default: edge_mask_reg_p6[487] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100001000,
	14'b1100100001001,
	14'b1100100001010,
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100011011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[488] <= 1'b1;
 		default: edge_mask_reg_p6[488] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100000,
	14'b1100100110000,
	14'b1100101000000,
	14'b1101100100000,
	14'b1101100110000,
	14'b1101101000000,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110101000000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000: edge_mask_reg_p6[489] <= 1'b1;
 		default: edge_mask_reg_p6[489] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1110100010000,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000: edge_mask_reg_p6[490] <= 1'b1;
 		default: edge_mask_reg_p6[490] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100000,
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011100000000,
	14'b10011100010000: edge_mask_reg_p6[491] <= 1'b1;
 		default: edge_mask_reg_p6[491] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100001,
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010001,
	14'b1111101010010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010001,
	14'b10010101010010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[492] <= 1'b1;
 		default: edge_mask_reg_p6[492] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100010,
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000001: edge_mask_reg_p6[493] <= 1'b1;
 		default: edge_mask_reg_p6[493] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100011,
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010011,
	14'b10010101010100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[494] <= 1'b1;
 		default: edge_mask_reg_p6[494] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100100,
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010100,
	14'b10010101010101,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000010,
	14'b10011101000011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001: edge_mask_reg_p6[495] <= 1'b1;
 		default: edge_mask_reg_p6[495] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100101,
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010101,
	14'b10010101010110,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000011,
	14'b10011101000100,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[496] <= 1'b1;
 		default: edge_mask_reg_p6[496] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100110,
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000100,
	14'b10011101000101,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[497] <= 1'b1;
 		default: edge_mask_reg_p6[497] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100100111,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[498] <= 1'b1;
 		default: edge_mask_reg_p6[498] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100011000,
	14'b1100100011001,
	14'b1100100011010,
	14'b1100100101000,
	14'b1100100101001,
	14'b1100100101010,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100011011,
	14'b1111100100000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000001,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[499] <= 1'b1;
 		default: edge_mask_reg_p6[499] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110000,
	14'b1100101000000,
	14'b1100101010000,
	14'b1101100110000,
	14'b1101101000000,
	14'b1101101010000,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000: edge_mask_reg_p6[500] <= 1'b1;
 		default: edge_mask_reg_p6[500] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110000,
	14'b1100100110001,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[501] <= 1'b1;
 		default: edge_mask_reg_p6[501] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110000,
	14'b1100100110001,
	14'b1100100110010,
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001: edge_mask_reg_p6[502] <= 1'b1;
 		default: edge_mask_reg_p6[502] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110001,
	14'b1100100110010,
	14'b1100100110011,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1110100100010,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100001,
	14'b1111101100010,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100001,
	14'b10000101100010,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100001,
	14'b10001101100010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100001,
	14'b10010101100010,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011101000000: edge_mask_reg_p6[503] <= 1'b1;
 		default: edge_mask_reg_p6[503] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110010,
	14'b1100100110011,
	14'b1100100110100,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1110100100011,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100010,
	14'b1111101100011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100010,
	14'b10000101100011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100010,
	14'b10001101100011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100010,
	14'b10010101100011,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10100100010000: edge_mask_reg_p6[504] <= 1'b1;
 		default: edge_mask_reg_p6[504] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110011,
	14'b1100100110100,
	14'b1100100110101,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100011,
	14'b1111101100100,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100011,
	14'b10000101100100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100011,
	14'b10001101100100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100011,
	14'b10010101100100,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[505] <= 1'b1;
 		default: edge_mask_reg_p6[505] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110100,
	14'b1100100110101,
	14'b1100100110110,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100100,
	14'b1111101100101,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100100,
	14'b10010101100101,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[506] <= 1'b1;
 		default: edge_mask_reg_p6[506] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110101,
	14'b1100100110110,
	14'b1100100110111,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100101,
	14'b10010101100110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[507] <= 1'b1;
 		default: edge_mask_reg_p6[507] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110110,
	14'b1100100110111,
	14'b1100100111000,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100110,
	14'b10010101100111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000: edge_mask_reg_p6[508] <= 1'b1;
 		default: edge_mask_reg_p6[508] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100110111,
	14'b1100100111000,
	14'b1100100111001,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100111,
	14'b10010101101000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000100,
	14'b10011101000101,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[509] <= 1'b1;
 		default: edge_mask_reg_p6[509] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100100111000,
	14'b1100100111001,
	14'b1100100111010,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100100000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100110000,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100101011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010100111011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[510] <= 1'b1;
 		default: edge_mask_reg_p6[510] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000000,
	14'b1100101010000,
	14'b1100101100000,
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101100000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000: edge_mask_reg_p6[511] <= 1'b1;
 		default: edge_mask_reg_p6[511] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[512] <= 1'b1;
 		default: edge_mask_reg_p6[512] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000000,
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001: edge_mask_reg_p6[513] <= 1'b1;
 		default: edge_mask_reg_p6[513] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000001,
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1110100110010,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110001,
	14'b1111101110010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110001,
	14'b10000101110010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110001,
	14'b10001101110010,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110001,
	14'b10010101110010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101010000: edge_mask_reg_p6[514] <= 1'b1;
 		default: edge_mask_reg_p6[514] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000010,
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1110100110011,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110010,
	14'b1111101110011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110010,
	14'b10000101110011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110010,
	14'b10001101110011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110010,
	14'b10010101110011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[515] <= 1'b1;
 		default: edge_mask_reg_p6[515] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000011,
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1110100110100,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110011,
	14'b1111101110100,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110011,
	14'b10000101110100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110011,
	14'b10001101110100,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110011,
	14'b10010101110100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000: edge_mask_reg_p6[516] <= 1'b1;
 		default: edge_mask_reg_p6[516] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000100,
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1110100110101,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110100,
	14'b1111101110101,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110100,
	14'b10000101110101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110100,
	14'b10001101110101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110100,
	14'b10010101110101,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[517] <= 1'b1;
 		default: edge_mask_reg_p6[517] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000101,
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1110100110110,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110101,
	14'b1111101110110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110101,
	14'b10000101110110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110101,
	14'b10001101110110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110101,
	14'b10010101110110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[518] <= 1'b1;
 		default: edge_mask_reg_p6[518] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000110,
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010100,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110110,
	14'b10010101110111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010011,
	14'b10011101010100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000: edge_mask_reg_p6[519] <= 1'b1;
 		default: edge_mask_reg_p6[519] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101000111,
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110111,
	14'b10010101111000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[520] <= 1'b1;
 		default: edge_mask_reg_p6[520] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101001000,
	14'b1100101001001,
	14'b1100101001010,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100110000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111100111011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010100111011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101111000,
	14'b10010101111001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[521] <= 1'b1;
 		default: edge_mask_reg_p6[521] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010000,
	14'b1100101100000,
	14'b1100101110000,
	14'b1101101010000,
	14'b1101101100000,
	14'b1101101110000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1110101110000,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000: edge_mask_reg_p6[522] <= 1'b1;
 		default: edge_mask_reg_p6[522] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011101000000: edge_mask_reg_p6[523] <= 1'b1;
 		default: edge_mask_reg_p6[523] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010000,
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000: edge_mask_reg_p6[524] <= 1'b1;
 		default: edge_mask_reg_p6[524] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010001,
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1110101000010,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000001,
	14'b1111110000010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000001,
	14'b10000110000010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000001,
	14'b10001110000010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000001,
	14'b10010110000010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101100000: edge_mask_reg_p6[525] <= 1'b1;
 		default: edge_mask_reg_p6[525] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010010,
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1110101000011,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000010,
	14'b1111110000011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000010,
	14'b10000110000011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000010,
	14'b10001110000011,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000010,
	14'b10010110000011,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10011101100001,
	14'b10100100000000,
	14'b10100100100000,
	14'b10100100110000: edge_mask_reg_p6[526] <= 1'b1;
 		default: edge_mask_reg_p6[526] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010011,
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1110101000100,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000011,
	14'b1111110000100,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000011,
	14'b10000110000100,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000011,
	14'b10001110000100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000011,
	14'b10010110000100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100001,
	14'b10011101100010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[527] <= 1'b1;
 		default: edge_mask_reg_p6[527] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010100,
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1110101000101,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000100,
	14'b1111110000101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000100,
	14'b10000110000101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000100,
	14'b10001110000101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000100,
	14'b10010110000101,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[528] <= 1'b1;
 		default: edge_mask_reg_p6[528] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010101,
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1110101000110,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000101,
	14'b1111110000110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000101,
	14'b10000110000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000101,
	14'b10001110000110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000101,
	14'b10010110000110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[529] <= 1'b1;
 		default: edge_mask_reg_p6[529] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010110,
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110101000111,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000110,
	14'b1111110000111,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000110,
	14'b10000110000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010000,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000110,
	14'b10001110000111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000110,
	14'b10010110000111,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100011,
	14'b10011101100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[530] <= 1'b1;
 		default: edge_mask_reg_p6[530] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101010111,
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010001,
	14'b1111100110000,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000000,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000111,
	14'b1111110001000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000111,
	14'b10000110001000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000111,
	14'b10001110001000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000111,
	14'b10010110001000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[531] <= 1'b1;
 		default: edge_mask_reg_p6[531] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101011000,
	14'b1100101011001,
	14'b1100101011010,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100110,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101001011,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110001000,
	14'b1111110001001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110001000,
	14'b10010110001001,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[532] <= 1'b1;
 		default: edge_mask_reg_p6[532] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100000,
	14'b1100101110000,
	14'b1100110000000,
	14'b1101101100000,
	14'b1101101110000,
	14'b1101110000000,
	14'b1110101100000,
	14'b1110101110000,
	14'b1110110000000,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010101000000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10011101000000,
	14'b10011101010000: edge_mask_reg_p6[533] <= 1'b1;
 		default: edge_mask_reg_p6[533] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110000001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101010000: edge_mask_reg_p6[534] <= 1'b1;
 		default: edge_mask_reg_p6[534] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100000,
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10001110010001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110010000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000: edge_mask_reg_p6[535] <= 1'b1;
 		default: edge_mask_reg_p6[535] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100001,
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1110101010010,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010001,
	14'b10000110010010,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010001,
	14'b10001110010010,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110010001,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101110000: edge_mask_reg_p6[536] <= 1'b1;
 		default: edge_mask_reg_p6[536] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100010,
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1110101010011,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010010,
	14'b1111110010011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010010,
	14'b10000110010011,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010010,
	14'b10001110010011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110010010,
	14'b10010110010011,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101110000,
	14'b10011101110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000: edge_mask_reg_p6[537] <= 1'b1;
 		default: edge_mask_reg_p6[537] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100011,
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1110101010100,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010011,
	14'b1111110010100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010011,
	14'b10000110010100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010011,
	14'b10001110010100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110010011,
	14'b10010110010100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110001,
	14'b10011101110010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[538] <= 1'b1;
 		default: edge_mask_reg_p6[538] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100100,
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1110101010101,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010100,
	14'b1111110010101,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010100,
	14'b10000110010101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010100,
	14'b10001110010101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110010100,
	14'b10010110010101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110010,
	14'b10011101110011,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[539] <= 1'b1;
 		default: edge_mask_reg_p6[539] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100101,
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1110101010110,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010101,
	14'b1111110010110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010101,
	14'b10000110010110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010101,
	14'b10001110010110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110010101,
	14'b10010110010110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[540] <= 1'b1;
 		default: edge_mask_reg_p6[540] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100110,
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101010111,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010110,
	14'b1111110010111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010110,
	14'b10000110010111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010110,
	14'b10001110010111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110010110,
	14'b10010110010111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100011,
	14'b10011101100100,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[541] <= 1'b1;
 		default: edge_mask_reg_p6[541] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101100111,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101011000,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000000,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010111,
	14'b1111110011000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010111,
	14'b10000110011000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010111,
	14'b10001110011000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110010111,
	14'b10010110011000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[542] <= 1'b1;
 		default: edge_mask_reg_p6[542] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100100000000,
	14'b1100101101000,
	14'b1100101101001,
	14'b1100101101010,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101011001,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101011011,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110011000,
	14'b1111110011001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110011000,
	14'b10000110011001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110011000,
	14'b10001110011001,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010101111011,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110011000,
	14'b10010110011001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010: edge_mask_reg_p6[543] <= 1'b1;
 		default: edge_mask_reg_p6[543] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110000,
	14'b1100110000000,
	14'b1100110010000,
	14'b1101101110000,
	14'b1101110000000,
	14'b1101110010000,
	14'b1110101110000,
	14'b1110110000000,
	14'b1110110010000,
	14'b1111101010000,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000101010000,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001101010000,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110010000,
	14'b10001110010001,
	14'b10010101010000,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110010000,
	14'b10011101010000,
	14'b10011101100000: edge_mask_reg_p6[544] <= 1'b1;
 		default: edge_mask_reg_p6[544] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110000,
	14'b1100101110001,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110010000,
	14'b1100110010001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110010000,
	14'b1101110010001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110100000,
	14'b10010101000000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110010000,
	14'b10010110010001,
	14'b10011101000000,
	14'b10011101010000,
	14'b10011101100000: edge_mask_reg_p6[545] <= 1'b1;
 		default: edge_mask_reg_p6[545] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110000,
	14'b1100101110001,
	14'b1100101110010,
	14'b1100110000000,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110010000,
	14'b1100110010001,
	14'b1100110010010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110010000,
	14'b1101110010001,
	14'b1101110010010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110100000,
	14'b1111110100001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10000110100001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110100000,
	14'b10001110100001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110010000,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110100000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10011101100001: edge_mask_reg_p6[546] <= 1'b1;
 		default: edge_mask_reg_p6[546] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110001,
	14'b1100101110010,
	14'b1100101110011,
	14'b1100110000001,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110010001,
	14'b1100110010010,
	14'b1100110010011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110010011,
	14'b1110101100010,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110100001,
	14'b1111110100010,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110100001,
	14'b10000110100010,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110100001,
	14'b10001110100010,
	14'b10010100010000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110010000,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110100001,
	14'b10011100010000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110000,
	14'b10100100010000,
	14'b10101100010000: edge_mask_reg_p6[547] <= 1'b1;
 		default: edge_mask_reg_p6[547] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110010,
	14'b1100101110011,
	14'b1100101110100,
	14'b1100110000010,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110010010,
	14'b1100110010011,
	14'b1100110010100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110010100,
	14'b1110101100011,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100000,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110100010,
	14'b1111110100011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110100010,
	14'b10000110100011,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110100010,
	14'b10001110100011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110000,
	14'b10011101110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[548] <= 1'b1;
 		default: edge_mask_reg_p6[548] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110011,
	14'b1100101110100,
	14'b1100101110101,
	14'b1100110000011,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110010011,
	14'b1100110010100,
	14'b1100110010101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110010101,
	14'b1110101100100,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100001,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110100011,
	14'b1111110100100,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110100011,
	14'b10000110100100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110100011,
	14'b10001110100100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110100011,
	14'b10010110100100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011110000001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[549] <= 1'b1;
 		default: edge_mask_reg_p6[549] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110100,
	14'b1100101110101,
	14'b1100101110110,
	14'b1100110000100,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110010100,
	14'b1100110010101,
	14'b1100110010110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110010110,
	14'b1110101100101,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110100100,
	14'b1111110100101,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110100100,
	14'b10000110100101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110100100,
	14'b10001110100101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110100100,
	14'b10010110100101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011110000010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[550] <= 1'b1;
 		default: edge_mask_reg_p6[550] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110101,
	14'b1100101110110,
	14'b1100101110111,
	14'b1100110000101,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110010101,
	14'b1100110010110,
	14'b1100110010111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110010111,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101100110,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110100101,
	14'b1111110100110,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110100101,
	14'b10000110100110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110100101,
	14'b10001110100110,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110100101,
	14'b10010110100110,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110010,
	14'b10011101110011,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[551] <= 1'b1;
 		default: edge_mask_reg_p6[551] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110110,
	14'b1100101110111,
	14'b1100101111000,
	14'b1100110000110,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110010110,
	14'b1100110010111,
	14'b1100110011000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110011000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101100111,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100001,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110100110,
	14'b1111110100111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110100110,
	14'b10000110100111,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110100110,
	14'b10001110100111,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110100110,
	14'b10010110100111,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[552] <= 1'b1;
 		default: edge_mask_reg_p6[552] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100101110111,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100110000111,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110010111,
	14'b1100110011000,
	14'b1100110011001,
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110011001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101101000,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100000,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110100111,
	14'b1111110101000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110100111,
	14'b10000110101000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110100111,
	14'b10001110101000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110011001,
	14'b10010110100111,
	14'b10010110101000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[553] <= 1'b1;
 		default: edge_mask_reg_p6[553] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100010000,
	14'b1100101111000,
	14'b1100101111001,
	14'b1100101111010,
	14'b1100110001000,
	14'b1100110001001,
	14'b1100110001010,
	14'b1100110011000,
	14'b1100110011001,
	14'b1100110011010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100010,
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110011000,
	14'b1101110011001,
	14'b1101110011010,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101101001,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110011010,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101101011,
	14'b1111101110000,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111101111011,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110001011,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110011010,
	14'b1111110101000,
	14'b1111110101001,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110000,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110001011,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110011010,
	14'b10000110101000,
	14'b10000110101001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110001011,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110011010,
	14'b10001110101000,
	14'b10001110101001,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010101111011,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110001011,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110011001,
	14'b10010110011010,
	14'b10010110101000,
	14'b10010110101001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010: edge_mask_reg_p6[554] <= 1'b1;
 		default: edge_mask_reg_p6[554] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100000,
	14'b1101001110000,
	14'b1101010000000,
	14'b1110001100000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1111001100000,
	14'b1111001110000,
	14'b1111010000000,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10010001100000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10011001100000,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000: edge_mask_reg_p6[555] <= 1'b1;
 		default: edge_mask_reg_p6[555] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b10000001010000,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10001001010000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010001010000,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10011001100000,
	14'b10011001100001,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10100010100000,
	14'b10100010110000: edge_mask_reg_p6[556] <= 1'b1;
 		default: edge_mask_reg_p6[556] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100000,
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1110001100000,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1111001100000,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b10000001010000,
	14'b10000001010001,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001010000,
	14'b10001001010001,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10010001010000,
	14'b10010001010001,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011001010000,
	14'b10011001100000,
	14'b10011001100001,
	14'b10011001100010,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10100010010000,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000: edge_mask_reg_p6[557] <= 1'b1;
 		default: edge_mask_reg_p6[557] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100001,
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1110001100001,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1111001100001,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b10000001010001,
	14'b10000001010010,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10001001010001,
	14'b10001001010010,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001010001,
	14'b10010001010010,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011001010001,
	14'b10011001100000,
	14'b10011001100001,
	14'b10011001100010,
	14'b10011001100011,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10100010000000,
	14'b10100010010000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000: edge_mask_reg_p6[558] <= 1'b1;
 		default: edge_mask_reg_p6[558] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100010,
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1110001100010,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1111001100010,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b10000001010010,
	14'b10000001010011,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110001,
	14'b10000010110010,
	14'b10001001010010,
	14'b10001001010011,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10010001010010,
	14'b10010001010011,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10011001010010,
	14'b10011001010011,
	14'b10011001100001,
	14'b10011001100010,
	14'b10011001100011,
	14'b10011001100100,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10100010000000,
	14'b10100010010000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10101011100000: edge_mask_reg_p6[559] <= 1'b1;
 		default: edge_mask_reg_p6[559] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100011,
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1110001100011,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1111001100011,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b10000001010011,
	14'b10000001010100,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110010,
	14'b10000010110011,
	14'b10001001010011,
	14'b10001001010100,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010001010011,
	14'b10010001010100,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011001010011,
	14'b10011001010100,
	14'b10011001100010,
	14'b10011001100011,
	14'b10011001100100,
	14'b10011001100101,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010000000,
	14'b10100010000001,
	14'b10100010010000,
	14'b10100010010001,
	14'b10100010010010,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[560] <= 1'b1;
 		default: edge_mask_reg_p6[560] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100100,
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1110001100100,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1111001100100,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b10000001010100,
	14'b10000001010101,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001010100,
	14'b10001001010101,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010001010100,
	14'b10010001010101,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011001010100,
	14'b10011001010101,
	14'b10011001100011,
	14'b10011001100100,
	14'b10011001100101,
	14'b10011001100110,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[561] <= 1'b1;
 		default: edge_mask_reg_p6[561] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100101,
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1110001100101,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1111001100101,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000001010101,
	14'b10000001010110,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001010101,
	14'b10001001010110,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010001010101,
	14'b10010001010110,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011001010101,
	14'b10011001010110,
	14'b10011001100100,
	14'b10011001100101,
	14'b10011001100110,
	14'b10011001100111,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101010110000,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[562] <= 1'b1;
 		default: edge_mask_reg_p6[562] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100110,
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1110001100110,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111001100110,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010110,
	14'b10000001010111,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001001010110,
	14'b10001001010111,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001010110,
	14'b10010001010111,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011001010110,
	14'b10011001010111,
	14'b10011001100101,
	14'b10011001100110,
	14'b10011001100111,
	14'b10011001101000,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10101011000000,
	14'b10101011010000: edge_mask_reg_p6[563] <= 1'b1;
 		default: edge_mask_reg_p6[563] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001100111,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110001100111,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111001100111,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010000,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b10000001010111,
	14'b10000001011000,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10001001010111,
	14'b10001001011000,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10010001010111,
	14'b10010001011000,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011001010111,
	14'b10011001011000,
	14'b10011001100110,
	14'b10011001100111,
	14'b10011001101000,
	14'b10011001101001,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011001111010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010001010,
	14'b10011010010000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000: edge_mask_reg_p6[564] <= 1'b1;
 		default: edge_mask_reg_p6[564] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011100000,
	14'b1100011100001,
	14'b1100011110000,
	14'b1100011110001,
	14'b1101001101000,
	14'b1101001101001,
	14'b1101001101010,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110001101000,
	14'b1110001101001,
	14'b1110001101010,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1111001101000,
	14'b1111001101001,
	14'b1111001101010,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001011000,
	14'b10000001011001,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001101010,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000001111011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001001011000,
	14'b10001001011001,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001101010,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001001111011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010001011000,
	14'b10010001011001,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001101010,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010001111011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010001011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10011001011000,
	14'b10011001011001,
	14'b10011001100111,
	14'b10011001101000,
	14'b10011001101001,
	14'b10011001101010,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011001111010,
	14'b10011001111011,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010001010,
	14'b10011010001011,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010011011,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000001,
	14'b10011011000010,
	14'b10100001101001,
	14'b10100001111001,
	14'b10100010001001: edge_mask_reg_p6[565] <= 1'b1;
 		default: edge_mask_reg_p6[565] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110000,
	14'b1101010000000,
	14'b1101010010000,
	14'b1110001110000,
	14'b1110010000000,
	14'b1110010010000,
	14'b1111001110000,
	14'b1111010000000,
	14'b1111010010000,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10010001110000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10011001110000,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000: edge_mask_reg_p6[566] <= 1'b1;
 		default: edge_mask_reg_p6[566] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110000,
	14'b1101001110001,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b10000001100000,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10001001100000,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001100000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10100010110000,
	14'b10100011000000: edge_mask_reg_p6[567] <= 1'b1;
 		default: edge_mask_reg_p6[567] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110000,
	14'b1101001110001,
	14'b1101001110010,
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1110001110000,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1111001110000,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b10000001100000,
	14'b10000001100001,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10001001100000,
	14'b10001001100001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010001100000,
	14'b10010001100001,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011001100000,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000: edge_mask_reg_p6[568] <= 1'b1;
 		default: edge_mask_reg_p6[568] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110001,
	14'b1101001110010,
	14'b1101001110011,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1110001110001,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1111001110001,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b10000001100001,
	14'b10000001100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10001001100001,
	14'b10001001100010,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10010001100001,
	14'b10010001100010,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011001100001,
	14'b10011001100010,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10100010010000,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001: edge_mask_reg_p6[569] <= 1'b1;
 		default: edge_mask_reg_p6[569] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110010,
	14'b1101001110011,
	14'b1101001110100,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1110001110010,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1111001110010,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b10000001100010,
	14'b10000001100011,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000001,
	14'b10001001100010,
	14'b10001001100011,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10010001100010,
	14'b10010001100011,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10011001100010,
	14'b10011001100011,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10100010010000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000: edge_mask_reg_p6[570] <= 1'b1;
 		default: edge_mask_reg_p6[570] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110011,
	14'b1101001110100,
	14'b1101001110101,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1110001110011,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1111001110011,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b10000001100011,
	14'b10000001100100,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000010,
	14'b10001001100011,
	14'b10001001100100,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10010001100011,
	14'b10010001100100,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011001100011,
	14'b10011001100100,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010010000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[571] <= 1'b1;
 		default: edge_mask_reg_p6[571] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110100,
	14'b1101001110101,
	14'b1101001110110,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1110001110100,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1111001110100,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b10000001100100,
	14'b10000001100101,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011110000,
	14'b10001001100100,
	14'b10001001100101,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011110000,
	14'b10010001100100,
	14'b10010001100101,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10011001100100,
	14'b10011001100101,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10100010010001,
	14'b10100010010010,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[572] <= 1'b1;
 		default: edge_mask_reg_p6[572] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110101,
	14'b1101001110110,
	14'b1101001110111,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1110001110101,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1111001110101,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111011110000,
	14'b10000001100101,
	14'b10000001100110,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011100000,
	14'b10000011110000,
	14'b10001001100101,
	14'b10001001100110,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010001100101,
	14'b10010001100110,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011001100101,
	14'b10011001100110,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000: edge_mask_reg_p6[573] <= 1'b1;
 		default: edge_mask_reg_p6[573] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110110,
	14'b1101001110111,
	14'b1101001111000,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1110001110110,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110011110000,
	14'b1111001110110,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000001100110,
	14'b10000001100111,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10001001100110,
	14'b10001001100111,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001100110,
	14'b10010001100111,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011001100110,
	14'b10011001100111,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[574] <= 1'b1;
 		default: edge_mask_reg_p6[574] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101001110111,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101011110000,
	14'b1110001110111,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1111001110111,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b10000001100111,
	14'b10000001101000,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001100111,
	14'b10001001101000,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001100111,
	14'b10010001101000,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011001100111,
	14'b10011001101000,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010001010,
	14'b10011010010000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000: edge_mask_reg_p6[575] <= 1'b1;
 		default: edge_mask_reg_p6[575] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1101001111000,
	14'b1101001111001,
	14'b1101001111010,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1110001111000,
	14'b1110001111001,
	14'b1110001111010,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1111001111000,
	14'b1111001111001,
	14'b1111001111010,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b10000001101000,
	14'b10000001101001,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000001111010,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010001011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001001101000,
	14'b10001001101001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010001011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001101000,
	14'b10010001101001,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010001011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011001101000,
	14'b10011001101001,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011001111010,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010001010,
	14'b10011010001011,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010011011,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010101011,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001: edge_mask_reg_p6[576] <= 1'b1;
 		default: edge_mask_reg_p6[576] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000000,
	14'b1101010010000,
	14'b1101010100000,
	14'b1110010000000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1111010000000,
	14'b1111010010000,
	14'b1111010100000,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10010010000000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10011010000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000: edge_mask_reg_p6[577] <= 1'b1;
 		default: edge_mask_reg_p6[577] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b10000001110000,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10001001110000,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10010001110000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10100011000000: edge_mask_reg_p6[578] <= 1'b1;
 		default: edge_mask_reg_p6[578] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000000,
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1110010000000,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1111010000000,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b10000001110000,
	14'b10000001110001,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001001110000,
	14'b10001001110001,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010001110000,
	14'b10010001110001,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011001110000,
	14'b10011001110001,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000: edge_mask_reg_p6[579] <= 1'b1;
 		default: edge_mask_reg_p6[579] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000001,
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1110010000001,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1111010000001,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b10000001110001,
	14'b10000001110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10001001110001,
	14'b10001001110010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010001110001,
	14'b10010001110010,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10011001110001,
	14'b10011001110010,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[580] <= 1'b1;
 		default: edge_mask_reg_p6[580] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000010,
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1110010000010,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1111010000010,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b10000001110010,
	14'b10000001110011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10001001110010,
	14'b10001001110011,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10010001110010,
	14'b10010001110011,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10011001110010,
	14'b10011001110011,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10100010010000,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001: edge_mask_reg_p6[581] <= 1'b1;
 		default: edge_mask_reg_p6[581] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000011,
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1110010000011,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1111010000011,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b10000001110011,
	14'b10000001110100,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10001001110011,
	14'b10001001110100,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10010001110011,
	14'b10010001110100,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10011001110011,
	14'b10011001110100,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010010001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[582] <= 1'b1;
 		default: edge_mask_reg_p6[582] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000100,
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1110010000100,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1111010000100,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b10000001110100,
	14'b10000001110101,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10001001110100,
	14'b10001001110101,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010001110100,
	14'b10010001110101,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011001110100,
	14'b10011001110101,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[583] <= 1'b1;
 		default: edge_mask_reg_p6[583] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000101,
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1110010000101,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1111010000101,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110110,
	14'b10000001110101,
	14'b10000001110110,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001001110101,
	14'b10001001110110,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10010001110101,
	14'b10010001110110,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011001110101,
	14'b10011001110110,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[584] <= 1'b1;
 		default: edge_mask_reg_p6[584] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000110,
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1110010000110,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1111010000110,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000001110110,
	14'b10000001110111,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010000,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001001110110,
	14'b10001001110111,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010001110110,
	14'b10010001110111,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011001110110,
	14'b10011001110111,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010100000,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000: edge_mask_reg_p6[585] <= 1'b1;
 		default: edge_mask_reg_p6[585] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010000111,
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1110010000111,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010000111,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010111000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001110111,
	14'b10000001111000,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001001110111,
	14'b10001001111000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010001110111,
	14'b10010001111000,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10011001110111,
	14'b10011001111000,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10101011000000,
	14'b10101011000001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[586] <= 1'b1;
 		default: edge_mask_reg_p6[586] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010001000,
	14'b1101010001001,
	14'b1101010001010,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010001000,
	14'b1110010001001,
	14'b1110010001010,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010001000,
	14'b1111010001001,
	14'b1111010001010,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000001111000,
	14'b10000001111001,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010011011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001001111000,
	14'b10001001111001,
	14'b10001001111010,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010011011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010001111000,
	14'b10010001111001,
	14'b10010001111010,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010011011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011001111000,
	14'b10011001111001,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010001010,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010011011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010101011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011010111011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[587] <= 1'b1;
 		default: edge_mask_reg_p6[587] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010000,
	14'b1101010100000,
	14'b1101010110000,
	14'b1110010010000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1111010010000,
	14'b1111010100000,
	14'b1111010110000,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001: edge_mask_reg_p6[588] <= 1'b1;
 		default: edge_mask_reg_p6[588] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b10000010000000,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10001010000000,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10010010000000,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10011010000000,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000: edge_mask_reg_p6[589] <= 1'b1;
 		default: edge_mask_reg_p6[589] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010000,
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1110010010000,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1111010010000,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b10000010000000,
	14'b10000010000001,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10001010000000,
	14'b10001010000001,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10010010000000,
	14'b10010010000001,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10011010000000,
	14'b10011010000001,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000: edge_mask_reg_p6[590] <= 1'b1;
 		default: edge_mask_reg_p6[590] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010001,
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1110010010001,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1111010010001,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b10000010000001,
	14'b10000010000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10001010000001,
	14'b10001010000010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10010010000001,
	14'b10010010000010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10011010000001,
	14'b10011010000010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10100010100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000: edge_mask_reg_p6[591] <= 1'b1;
 		default: edge_mask_reg_p6[591] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010010,
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1110010010010,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1111010010010,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b10000010000010,
	14'b10000010000011,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10001010000010,
	14'b10001010000011,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010000010,
	14'b10010010000011,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10011010000010,
	14'b10011010000011,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[592] <= 1'b1;
 		default: edge_mask_reg_p6[592] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010011,
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1110010010011,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1111010010011,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000100,
	14'b10000010000011,
	14'b10000010000100,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10001010000011,
	14'b10001010000100,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010000011,
	14'b10010010000100,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10011010000011,
	14'b10011010000100,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10100010100000,
	14'b10100010100001,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[593] <= 1'b1;
 		default: edge_mask_reg_p6[593] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010100,
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1110010010100,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1111010010100,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000101,
	14'b10000010000100,
	14'b10000010000101,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10001010000100,
	14'b10001010000101,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010000100,
	14'b10010010000101,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010100000000,
	14'b10011010000100,
	14'b10011010000101,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100010100001,
	14'b10100010100010,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[594] <= 1'b1;
 		default: edge_mask_reg_p6[594] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010101,
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1110010010101,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1111010010101,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000110,
	14'b10000010000101,
	14'b10000010000110,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000100000000,
	14'b10001010000101,
	14'b10001010000110,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001100000000,
	14'b10010010000101,
	14'b10010010000110,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10011010000101,
	14'b10011010000110,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10100010100010,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10110011100000: edge_mask_reg_p6[595] <= 1'b1;
 		default: edge_mask_reg_p6[595] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010110,
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1110010010110,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1111010010110,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000111,
	14'b1111011110000,
	14'b1111100000000,
	14'b10000010000110,
	14'b10000010000111,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10001010000110,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010000110,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010000110,
	14'b10011010000111,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011000000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[596] <= 1'b1;
 		default: edge_mask_reg_p6[596] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010010111,
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1110010010111,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111010010111,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011001000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b10000010000111,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010000111,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100000,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010000111,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010000111,
	14'b10011010001000,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010100000,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001: edge_mask_reg_p6[597] <= 1'b1;
 		default: edge_mask_reg_p6[597] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010011000,
	14'b1101010011001,
	14'b1101010011010,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110010011000,
	14'b1110010011001,
	14'b1110010011010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111010011000,
	14'b1111010011001,
	14'b1111010011010,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011001001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b10000010001000,
	14'b10000010001001,
	14'b10000010001010,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010101011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010001000,
	14'b10001010001001,
	14'b10001010001010,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010101011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010001000,
	14'b10010010001001,
	14'b10010010001010,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010101011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011001011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010001000,
	14'b10011010001001,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010101011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011010111011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011001011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000: edge_mask_reg_p6[598] <= 1'b1;
 		default: edge_mask_reg_p6[598] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100000,
	14'b1101010110000,
	14'b1101011000000,
	14'b1110010100000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1111010100000,
	14'b1111010110000,
	14'b1111011000000,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001: edge_mask_reg_p6[599] <= 1'b1;
 		default: edge_mask_reg_p6[599] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b10000010010000,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10001010010000,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10010010010000,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10011010010000,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000: edge_mask_reg_p6[600] <= 1'b1;
 		default: edge_mask_reg_p6[600] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100000,
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1110010100000,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1111010100000,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b10000010010000,
	14'b10000010010001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010010000,
	14'b10001010010001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10010010010000,
	14'b10010010010001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10011010010000,
	14'b10011010010001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10100011010000,
	14'b10100011100000: edge_mask_reg_p6[601] <= 1'b1;
 		default: edge_mask_reg_p6[601] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100001,
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1110010100001,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1111010100001,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b10000010010001,
	14'b10000010010010,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10001010010001,
	14'b10001010010010,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010010010001,
	14'b10010010010010,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011010010001,
	14'b10011010010010,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001: edge_mask_reg_p6[602] <= 1'b1;
 		default: edge_mask_reg_p6[602] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100010,
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1110010100010,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1111010100010,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010011,
	14'b10000010010010,
	14'b10000010010011,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10001010010010,
	14'b10001010010011,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10010010010010,
	14'b10010010010011,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10011010010010,
	14'b10011010010011,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000: edge_mask_reg_p6[603] <= 1'b1;
 		default: edge_mask_reg_p6[603] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100011,
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1110010100011,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1111010100011,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010100,
	14'b10000010010011,
	14'b10000010010100,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10001010010011,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10010010010011,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10011010010011,
	14'b10011010010100,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10100010110000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000: edge_mask_reg_p6[604] <= 1'b1;
 		default: edge_mask_reg_p6[604] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100100,
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1110010100100,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1111010100100,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010101,
	14'b10000010010100,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10001010010100,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10010010010100,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10011010010100,
	14'b10011010010101,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10100010110001,
	14'b10100010110010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[605] <= 1'b1;
 		default: edge_mask_reg_p6[605] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100101,
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1110010100101,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1111010100101,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010110,
	14'b10000010010101,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10001010010101,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010010101,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011010010101,
	14'b10011010010110,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100010110010,
	14'b10100010110011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011010100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[606] <= 1'b1;
 		default: edge_mask_reg_p6[606] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100110,
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1110010100110,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1111010100110,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010111,
	14'b10000010010110,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010010110,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10010010010110,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010010110,
	14'b10011010010111,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[607] <= 1'b1;
 		default: edge_mask_reg_p6[607] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010100111,
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1110010100111,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1111010100111,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011011000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010010111,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110000,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10001010010111,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010010010111,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011010010111,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[608] <= 1'b1;
 		default: edge_mask_reg_p6[608] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010101000,
	14'b1101010101001,
	14'b1101010101010,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1110010101000,
	14'b1110010101001,
	14'b1110010101010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010101000,
	14'b1111010101001,
	14'b1111010101010,
	14'b1111010110000,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011011001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010011000,
	14'b10000010011001,
	14'b10000010011010,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000010111011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010011000,
	14'b10001010011001,
	14'b10001010011010,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001010111011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010010011000,
	14'b10010010011001,
	14'b10010010011010,
	14'b10010010100000,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010010111011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011001011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011011011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011010011000,
	14'b10011010011001,
	14'b10011010011010,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011010111011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011001011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011011011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001: edge_mask_reg_p6[609] <= 1'b1;
 		default: edge_mask_reg_p6[609] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110000,
	14'b1101011000000,
	14'b1101011010000,
	14'b1110010110000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1111010110000,
	14'b1111011000000,
	14'b1111011010000,
	14'b10000010110000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10001010110000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10010010110000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001: edge_mask_reg_p6[610] <= 1'b1;
 		default: edge_mask_reg_p6[610] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110000,
	14'b1101010110001,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b10000010100000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10001010100000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10010010100000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10011010100000,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000: edge_mask_reg_p6[611] <= 1'b1;
 		default: edge_mask_reg_p6[611] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110000,
	14'b1101010110001,
	14'b1101010110010,
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1110010110000,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1111010110000,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100001,
	14'b10000010100000,
	14'b10000010100001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001010100000,
	14'b10001010100001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010010100000,
	14'b10010010100001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10011010100000,
	14'b10011010100001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001: edge_mask_reg_p6[612] <= 1'b1;
 		default: edge_mask_reg_p6[612] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110001,
	14'b1101010110010,
	14'b1101010110011,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1110010110001,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1111010110001,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100010,
	14'b10000010100001,
	14'b10000010100010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10001010100001,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10010010100001,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10011010100001,
	14'b10011010100010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001: edge_mask_reg_p6[613] <= 1'b1;
 		default: edge_mask_reg_p6[613] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110010,
	14'b1101010110011,
	14'b1101010110100,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1110010110010,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1111010110010,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100011,
	14'b10000010100010,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10001010100010,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10010010100010,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10011010100010,
	14'b10011010100011,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010: edge_mask_reg_p6[614] <= 1'b1;
 		default: edge_mask_reg_p6[614] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110011,
	14'b1101010110100,
	14'b1101010110101,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1110010110011,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1111010110011,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100100,
	14'b10000010100011,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10001010100011,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10010010100011,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10011010100011,
	14'b10011010100100,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10100010110001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010: edge_mask_reg_p6[615] <= 1'b1;
 		default: edge_mask_reg_p6[615] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110100,
	14'b1101010110101,
	14'b1101010110110,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1110010110100,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1111010110100,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100101,
	14'b10000010100100,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010010,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10001010100100,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10010010100100,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10011010100100,
	14'b10011010100101,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000: edge_mask_reg_p6[616] <= 1'b1;
 		default: edge_mask_reg_p6[616] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110101,
	14'b1101010110110,
	14'b1101010110111,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1110010110101,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1111010110101,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100110,
	14'b10000010100101,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100010000,
	14'b10011010100101,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100010000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100010000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[617] <= 1'b1;
 		default: edge_mask_reg_p6[617] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110110,
	14'b1101010110111,
	14'b1101010111000,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1110010110110,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1111010110110,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100111,
	14'b10000010100110,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000000,
	14'b10000100010000,
	14'b10001010100101,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100010000,
	14'b10010010100101,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010110000,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011010100110,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010110000,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011010100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[618] <= 1'b1;
 		default: edge_mask_reg_p6[618] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010110111,
	14'b1101010111000,
	14'b1101010111001,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1110010110111,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1111010110111,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011101000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010100111,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001010100110,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010110000,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10010010100110,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010100111,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011010001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[619] <= 1'b1;
 		default: edge_mask_reg_p6[619] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101010111000,
	14'b1101010111001,
	14'b1101010111010,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1110010111000,
	14'b1110010111001,
	14'b1110010111010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111010111000,
	14'b1111010111001,
	14'b1111010111010,
	14'b1111011000000,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011101001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010101000,
	14'b10000010101001,
	14'b10000010101010,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011001011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010100111,
	14'b10001010101000,
	14'b10001010101001,
	14'b10001010101010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011001011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010010100111,
	14'b10010010101000,
	14'b10010010101001,
	14'b10010010101010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011001011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011011011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011101011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010101000,
	14'b10011010101001,
	14'b10011010101010,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011011011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100010110000,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[620] <= 1'b1;
 		default: edge_mask_reg_p6[620] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000000,
	14'b1101011010000,
	14'b1101011100000,
	14'b1110011000000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011100000,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001: edge_mask_reg_p6[621] <= 1'b1;
 		default: edge_mask_reg_p6[621] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10011010110000,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000: edge_mask_reg_p6[622] <= 1'b1;
 		default: edge_mask_reg_p6[622] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000000,
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1110011000000,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1111011000000,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110001,
	14'b10000010110000,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011010110000,
	14'b10011010110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001: edge_mask_reg_p6[623] <= 1'b1;
 		default: edge_mask_reg_p6[623] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000001,
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1110011000001,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1111011000001,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110010,
	14'b10000010110001,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10011010110001,
	14'b10011010110010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[624] <= 1'b1;
 		default: edge_mask_reg_p6[624] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000010,
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1110011000010,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1111011000010,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110011,
	14'b10000010110010,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10001010110001,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10010010110001,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10011010110010,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001: edge_mask_reg_p6[625] <= 1'b1;
 		default: edge_mask_reg_p6[625] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000011,
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1110011000011,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1111011000011,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110100,
	14'b10000010110011,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10001010110010,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10010010110010,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10011010110011,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010: edge_mask_reg_p6[626] <= 1'b1;
 		default: edge_mask_reg_p6[626] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000100,
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1110011000100,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1111011000100,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110101,
	14'b10000010110100,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10001010110011,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10010010110011,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10011010110100,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10100011000001,
	14'b10100011000010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011: edge_mask_reg_p6[627] <= 1'b1;
 		default: edge_mask_reg_p6[627] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000101,
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1110011000101,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1111011000101,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110110,
	14'b10000010110101,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10001010110100,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10010010110100,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10011010110101,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10100011000010,
	14'b10100011000011,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000: edge_mask_reg_p6[628] <= 1'b1;
 		default: edge_mask_reg_p6[628] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000110,
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1110011000110,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1111011000110,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110111,
	14'b10000010110110,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10001010110101,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10010010110101,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010011000000,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10011010110110,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011011000000,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011010100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011100000,
	14'b10110011110000: edge_mask_reg_p6[629] <= 1'b1;
 		default: edge_mask_reg_p6[629] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011000111,
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1110011000111,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1111011000111,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011111000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000010110111,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000011000000,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000000,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10001010110110,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10010010110110,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011010110111,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[630] <= 1'b1;
 		default: edge_mask_reg_p6[630] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011001000,
	14'b1101011001001,
	14'b1101011001010,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1110011001000,
	14'b1110011001001,
	14'b1110011001010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110100000000,
	14'b1110100010000,
	14'b1111011000000,
	14'b1111011001000,
	14'b1111011001001,
	14'b1111011001010,
	14'b1111011010000,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011111001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000010111000,
	14'b10000010111001,
	14'b10000010111010,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011011011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001010110000,
	14'b10001010110001,
	14'b10001010110111,
	14'b10001010111000,
	14'b10001010111001,
	14'b10001010111010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010010110000,
	14'b10010010110001,
	14'b10010010110111,
	14'b10010010111000,
	14'b10010010111001,
	14'b10010010111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011011011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011101011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011010110000,
	14'b10011010111000,
	14'b10011010111001,
	14'b10011010111010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011101011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011011111010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001: edge_mask_reg_p6[631] <= 1'b1;
 		default: edge_mask_reg_p6[631] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010000,
	14'b1101011100000,
	14'b1101011110000,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011110000,
	14'b10000011000000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10001011000000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000: edge_mask_reg_p6[632] <= 1'b1;
 		default: edge_mask_reg_p6[632] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001: edge_mask_reg_p6[633] <= 1'b1;
 		default: edge_mask_reg_p6[633] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010000,
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1110011010000,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1111011010000,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000001,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010: edge_mask_reg_p6[634] <= 1'b1;
 		default: edge_mask_reg_p6[634] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010001,
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1110011010001,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1111011010001,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000010,
	14'b10000011000001,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000: edge_mask_reg_p6[635] <= 1'b1;
 		default: edge_mask_reg_p6[635] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010010,
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1110011010010,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1111011010010,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000011,
	14'b10000011000010,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10011011000010,
	14'b10011011000011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000: edge_mask_reg_p6[636] <= 1'b1;
 		default: edge_mask_reg_p6[636] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010011,
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1110011010011,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1111011010011,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000100,
	14'b10000011000011,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10001011000010,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10010011000010,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10011011000011,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010: edge_mask_reg_p6[637] <= 1'b1;
 		default: edge_mask_reg_p6[637] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010100,
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1110011010100,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1111011010100,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000101,
	14'b1111100000110,
	14'b10000011000100,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10001011000011,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10010011000011,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10100011010001,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011: edge_mask_reg_p6[638] <= 1'b1;
 		default: edge_mask_reg_p6[638] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010101,
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1110011010101,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1111011010101,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000110,
	14'b1111100000111,
	14'b10000011000101,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10001011000100,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10010011000100,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10011011000100,
	14'b10011011000101,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10100011010000,
	14'b10100011010010,
	14'b10100011010011,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000: edge_mask_reg_p6[639] <= 1'b1;
 		default: edge_mask_reg_p6[639] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010110,
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1110011010110,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1111011010110,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000111,
	14'b1111100001000,
	14'b10000011000110,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10001011000101,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10010011000000,
	14'b10010011000101,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10011011000000,
	14'b10011011000110,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010011,
	14'b10100011010100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100100000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[640] <= 1'b1;
 		default: edge_mask_reg_p6[640] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011010111,
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1110011010111,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1111011010111,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100001000,
	14'b1111100001001,
	14'b10000011000000,
	14'b10000011000111,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011010000,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000110,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000110,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000111,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[641] <= 1'b1;
 		default: edge_mask_reg_p6[641] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011011000,
	14'b1101011011001,
	14'b1101011011010,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1110011011000,
	14'b1110011011001,
	14'b1110011011010,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100010000,
	14'b1111011000000,
	14'b1111011010000,
	14'b1111011011000,
	14'b1111011011001,
	14'b1111011011010,
	14'b1111011100000,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100000000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100100000,
	14'b10000011000000,
	14'b10000011000001,
	14'b10000011001000,
	14'b10000011001001,
	14'b10000011001010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011000010,
	14'b10001011000111,
	14'b10001011001000,
	14'b10001011001001,
	14'b10001011001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011011011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011000010,
	14'b10010011000111,
	14'b10010011001000,
	14'b10010011001001,
	14'b10010011001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011011011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011101011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010011111011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011000010,
	14'b10011011001000,
	14'b10011011001001,
	14'b10011011001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011011111010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10100011000000,
	14'b10100011000001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011100000,
	14'b10101011100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[642] <= 1'b1;
 		default: edge_mask_reg_p6[642] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100000,
	14'b1101011110000,
	14'b1101100000000,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100100000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000: edge_mask_reg_p6[643] <= 1'b1;
 		default: edge_mask_reg_p6[643] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001: edge_mask_reg_p6[644] <= 1'b1;
 		default: edge_mask_reg_p6[644] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100000,
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1110011100000,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010001,
	14'b1111100010010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010: edge_mask_reg_p6[645] <= 1'b1;
 		default: edge_mask_reg_p6[645] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100001,
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1110011100001,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1111011100001,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b10000011010001,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000: edge_mask_reg_p6[646] <= 1'b1;
 		default: edge_mask_reg_p6[646] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100010,
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1110011100010,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1111011100010,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b10000011010010,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001: edge_mask_reg_p6[647] <= 1'b1;
 		default: edge_mask_reg_p6[647] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100011,
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1110011100011,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1111011100011,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b10000011010011,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10001011010010,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10010011010010,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10011011010010,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010: edge_mask_reg_p6[648] <= 1'b1;
 		default: edge_mask_reg_p6[648] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100100,
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1110011100100,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1111011100100,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b10000011010100,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10001011010011,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10010011010011,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10011011010011,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011: edge_mask_reg_p6[649] <= 1'b1;
 		default: edge_mask_reg_p6[649] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100101,
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1110011100101,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1111011100101,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010110,
	14'b1111100010111,
	14'b10000011010101,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10001011010100,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10010011010100,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10011011010100,
	14'b10011011010101,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011: edge_mask_reg_p6[650] <= 1'b1;
 		default: edge_mask_reg_p6[650] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100110,
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1110011100110,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1111011100110,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010111,
	14'b1111100011000,
	14'b10000011010110,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10001011010000,
	14'b10001011010101,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10010011010000,
	14'b10010011010101,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10011011010000,
	14'b10011011010110,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011100011,
	14'b10100011100100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110011110000,
	14'b10110100000000: edge_mask_reg_p6[651] <= 1'b1;
 		default: edge_mask_reg_p6[651] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011100111,
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1110011100111,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1111011100111,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100011000,
	14'b1111100011001,
	14'b10000011010000,
	14'b10000011010111,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011100000,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010110,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010110,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010111,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10100011000000,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[652] <= 1'b1;
 		default: edge_mask_reg_p6[652] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011101000,
	14'b1101011101001,
	14'b1101011101010,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1110011101000,
	14'b1110011101001,
	14'b1110011101010,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011101000,
	14'b1111011101001,
	14'b1111011101010,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011011000,
	14'b10000011011001,
	14'b10000011011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011101011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10001011000000,
	14'b10001011000001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011010111,
	14'b10001011011000,
	14'b10001011011001,
	14'b10001011011010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011101011,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100001011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011010111,
	14'b10010011011000,
	14'b10010011011001,
	14'b10010011011010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011101011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010011111011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100001011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011000000,
	14'b10011011000001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011011000,
	14'b10011011011001,
	14'b10011011011010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011011111010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001: edge_mask_reg_p6[653] <= 1'b1;
 		default: edge_mask_reg_p6[653] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000000,
	14'b1101100010000,
	14'b1101100100000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110100100000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111100100000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000: edge_mask_reg_p6[654] <= 1'b1;
 		default: edge_mask_reg_p6[654] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001: edge_mask_reg_p6[655] <= 1'b1;
 		default: edge_mask_reg_p6[655] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110000,
	14'b1101011110001,
	14'b1101011110010,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010: edge_mask_reg_p6[656] <= 1'b1;
 		default: edge_mask_reg_p6[656] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110001,
	14'b1101011110010,
	14'b1101011110011,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1110011110001,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[657] <= 1'b1;
 		default: edge_mask_reg_p6[657] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110010,
	14'b1101011110011,
	14'b1101011110100,
	14'b1101100000010,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1110011110010,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1111011110010,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001: edge_mask_reg_p6[658] <= 1'b1;
 		default: edge_mask_reg_p6[658] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110011,
	14'b1101011110100,
	14'b1101011110101,
	14'b1101100000011,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1110011110011,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110100000011,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1111011110011,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b10000011100010,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010: edge_mask_reg_p6[659] <= 1'b1;
 		default: edge_mask_reg_p6[659] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110100,
	14'b1101011110101,
	14'b1101011110110,
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1110011110100,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1111011110100,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10011011100000,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011: edge_mask_reg_p6[660] <= 1'b1;
 		default: edge_mask_reg_p6[660] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110101,
	14'b1101011110110,
	14'b1101011110111,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1110011110101,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1111011110101,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b10000011100011,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10010011100000,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100011,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100010,
	14'b10100100100011: edge_mask_reg_p6[661] <= 1'b1;
 		default: edge_mask_reg_p6[661] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110110,
	14'b1101011110111,
	14'b1101011111000,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1110011110110,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1111011110110,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b10000011100100,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011100011,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100011,
	14'b10010011100100,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100100,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100110000,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10100100100011,
	14'b10100100100100,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10110011110000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[662] <= 1'b1;
 		default: edge_mask_reg_p6[662] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110111,
	14'b1101011111000,
	14'b1101011111001,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1110011110111,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1111011110111,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100100,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10010011000000,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100101,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10011011000000,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100101,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000: edge_mask_reg_p6[663] <= 1'b1;
 		default: edge_mask_reg_p6[663] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011111000,
	14'b1101011111001,
	14'b1101011111010,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1110011010000,
	14'b1110011100000,
	14'b1110011111000,
	14'b1110011111001,
	14'b1110011111010,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011111000,
	14'b1111011111001,
	14'b1111011111010,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100010000,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100101,
	14'b10000011100110,
	14'b10000011100111,
	14'b10000011101000,
	14'b10000011101001,
	14'b10000011101010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000011111011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100001011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011010010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011100101,
	14'b10001011100110,
	14'b10001011100111,
	14'b10001011101000,
	14'b10001011101001,
	14'b10001011101010,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001011111011,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100001011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10010011000000,
	14'b10010011000001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011100110,
	14'b10010011100111,
	14'b10010011101000,
	14'b10010011101001,
	14'b10010011101010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010011111011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100001011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100011011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011010010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011100110,
	14'b10011011100111,
	14'b10011011101000,
	14'b10011011101001,
	14'b10011011101010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011011111010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100001011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[664] <= 1'b1;
 		default: edge_mask_reg_p6[664] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010000,
	14'b1101100100000,
	14'b1101100110000,
	14'b1110100010000,
	14'b1110100100000,
	14'b1110100110000,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100110000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000: edge_mask_reg_p6[665] <= 1'b1;
 		default: edge_mask_reg_p6[665] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000: edge_mask_reg_p6[666] <= 1'b1;
 		default: edge_mask_reg_p6[666] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001: edge_mask_reg_p6[667] <= 1'b1;
 		default: edge_mask_reg_p6[667] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000001,
	14'b10011101000010,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[668] <= 1'b1;
 		default: edge_mask_reg_p6[668] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[669] <= 1'b1;
 		default: edge_mask_reg_p6[669] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100010011,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1111100000011,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[670] <= 1'b1;
 		default: edge_mask_reg_p6[670] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000100,
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100010100,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1110100000100,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100010100,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1111100000100,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010010,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110010: edge_mask_reg_p6[671] <= 1'b1;
 		default: edge_mask_reg_p6[671] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000101,
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100010101,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1110100000101,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100010101,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1111100000101,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b10000011110011,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100011110100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110011: edge_mask_reg_p6[672] <= 1'b1;
 		default: edge_mask_reg_p6[672] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000110,
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100010110,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1110100000110,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100010110,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1111100000110,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10001011010000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100110000,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100011110011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100100100,
	14'b10100100110000,
	14'b10101011010000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[673] <= 1'b1;
 		default: edge_mask_reg_p6[673] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000111,
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100010111,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1110100000111,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100010111,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100000111,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b10000011010000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110100,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011101000000,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101011110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000: edge_mask_reg_p6[674] <= 1'b1;
 		default: edge_mask_reg_p6[674] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100001000,
	14'b1101100001001,
	14'b1101100001010,
	14'b1101100011000,
	14'b1101100011001,
	14'b1101100011010,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100001000,
	14'b1110100001001,
	14'b1110100001010,
	14'b1110100011000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1111011010000,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100001000,
	14'b1111100001001,
	14'b1111100001010,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b10000011010000,
	14'b10000011010001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000011110101,
	14'b10000011110110,
	14'b10000011110111,
	14'b10000011111000,
	14'b10000011111001,
	14'b10000011111010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001011110100,
	14'b10001011110101,
	14'b10001011110110,
	14'b10001011110111,
	14'b10001011111000,
	14'b10001011111001,
	14'b10001011111010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100001011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011010010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010011110100,
	14'b10010011110101,
	14'b10010011110110,
	14'b10010011110111,
	14'b10010011111000,
	14'b10010011111001,
	14'b10010011111010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100001011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100011011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011011110100,
	14'b10011011110101,
	14'b10011011110110,
	14'b10011011110111,
	14'b10011011111000,
	14'b10011011111001,
	14'b10011011111010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100011011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10100011010000,
	14'b10100011010001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[675] <= 1'b1;
 		default: edge_mask_reg_p6[675] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100000,
	14'b1101100110000,
	14'b1101101000000,
	14'b1110100100000,
	14'b1110100110000,
	14'b1110101000000,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111101000000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000: edge_mask_reg_p6[676] <= 1'b1;
 		default: edge_mask_reg_p6[676] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1111100010000,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000: edge_mask_reg_p6[677] <= 1'b1;
 		default: edge_mask_reg_p6[677] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10100100000000: edge_mask_reg_p6[678] <= 1'b1;
 		default: edge_mask_reg_p6[678] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010001,
	14'b10000101010010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010001,
	14'b10011101010010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000: edge_mask_reg_p6[679] <= 1'b1;
 		default: edge_mask_reg_p6[679] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100000,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010010,
	14'b10011101010011,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[680] <= 1'b1;
 		default: edge_mask_reg_p6[680] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100011,
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1111100010100,
	14'b1111100010101,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100001,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010011,
	14'b10011101010100,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[681] <= 1'b1;
 		default: edge_mask_reg_p6[681] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100100,
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1110100100100,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1111100010101,
	14'b1111100010110,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010100,
	14'b10011101010101,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011: edge_mask_reg_p6[682] <= 1'b1;
 		default: edge_mask_reg_p6[682] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100101,
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1110100100101,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1111100010110,
	14'b1111100010111,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[683] <= 1'b1;
 		default: edge_mask_reg_p6[683] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100110,
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1110100100110,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1111100010111,
	14'b1111100011000,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10100011010000,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100000011,
	14'b10100100000100,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100100100,
	14'b10100100110000,
	14'b10100100110011,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110100000000,
	14'b10110100010000: edge_mask_reg_p6[684] <= 1'b1;
 		default: edge_mask_reg_p6[684] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100100111,
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1110100100111,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100011000,
	14'b1111100011001,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100010000,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10010011010000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011101000000,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[685] <= 1'b1;
 		default: edge_mask_reg_p6[685] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100101000,
	14'b1101100101001,
	14'b1101100101010,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100011001,
	14'b1110100011010,
	14'b1110100101000,
	14'b1110100101001,
	14'b1110100101010,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100011001,
	14'b1111100011010,
	14'b1111100100000,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100000100,
	14'b10000100000101,
	14'b10000100000110,
	14'b10000100000111,
	14'b10000100001000,
	14'b10000100001001,
	14'b10000100001010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100011011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10001011010000,
	14'b10001011010001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011100011,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100000101,
	14'b10001100000110,
	14'b10001100000111,
	14'b10001100001000,
	14'b10001100001001,
	14'b10001100001010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100011011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10010011010000,
	14'b10010011010001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011100011,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100000101,
	14'b10010100000110,
	14'b10010100000111,
	14'b10010100001000,
	14'b10010100001001,
	14'b10010100001010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100011011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010100111011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10011011010000,
	14'b10011011010001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011100011,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100000100,
	14'b10011100000101,
	14'b10011100000110,
	14'b10011100000111,
	14'b10011100001000,
	14'b10011100001001,
	14'b10011100001010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100101011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011100010,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001: edge_mask_reg_p6[686] <= 1'b1;
 		default: edge_mask_reg_p6[686] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110000,
	14'b1101101000000,
	14'b1101101010000,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101010000,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000: edge_mask_reg_p6[687] <= 1'b1;
 		default: edge_mask_reg_p6[687] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110000,
	14'b1101100110001,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1111100100000,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000: edge_mask_reg_p6[688] <= 1'b1;
 		default: edge_mask_reg_p6[688] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10100100010000,
	14'b10100100100000: edge_mask_reg_p6[689] <= 1'b1;
 		default: edge_mask_reg_p6[689] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1111100100010,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100001,
	14'b10000101100010,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100001,
	14'b10001101100010,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100001,
	14'b10010101100010,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100001,
	14'b10011101100010,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100101000000: edge_mask_reg_p6[690] <= 1'b1;
 		default: edge_mask_reg_p6[690] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110010,
	14'b1101100110011,
	14'b1101100110100,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1111100100011,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100010,
	14'b10000101100011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100010,
	14'b10001101100011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100010,
	14'b10010101100011,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100010,
	14'b10011101100011,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[691] <= 1'b1;
 		default: edge_mask_reg_p6[691] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110011,
	14'b1101100110100,
	14'b1101100110101,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1111100100100,
	14'b1111100100101,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100011,
	14'b10000101100100,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100011,
	14'b10011101100100,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010: edge_mask_reg_p6[692] <= 1'b1;
 		default: edge_mask_reg_p6[692] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110100,
	14'b1101100110101,
	14'b1101100110110,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1110100110100,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1111100100101,
	14'b1111100100110,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101100100,
	14'b10011101100101,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000001,
	14'b10100101000010: edge_mask_reg_p6[693] <= 1'b1;
 		default: edge_mask_reg_p6[693] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110101,
	14'b1101100110110,
	14'b1101100110111,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1110100110101,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1111100100110,
	14'b1111100100111,
	14'b1111100110101,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101100101,
	14'b10011101100110,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100010100,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100100100,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000010,
	14'b10100101000011,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[694] <= 1'b1;
 		default: edge_mask_reg_p6[694] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110110,
	14'b1101100110111,
	14'b1101100111000,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1110100110110,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1111100100111,
	14'b1111100101000,
	14'b1111100110110,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10011011010000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011101000000,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101100110,
	14'b10011101100111,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100010011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10110100010000: edge_mask_reg_p6[695] <= 1'b1;
 		default: edge_mask_reg_p6[695] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100110111,
	14'b1101100111000,
	14'b1101100111001,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1110100110111,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111100101000,
	14'b1111100101001,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100100000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10100011100000,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[696] <= 1'b1;
 		default: edge_mask_reg_p6[696] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100111000,
	14'b1101100111001,
	14'b1101100111010,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110100111000,
	14'b1110100111001,
	14'b1110100111010,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1111011100000,
	14'b1111011100001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000001,
	14'b1111100100000,
	14'b1111100101001,
	14'b1111100101010,
	14'b1111100110000,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b10000011100000,
	14'b10000011100001,
	14'b10000011100010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100010101,
	14'b10000100010110,
	14'b10000100010111,
	14'b10000100011000,
	14'b10000100011001,
	14'b10000100011010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100101011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100010101,
	14'b10001100010110,
	14'b10001100010111,
	14'b10001100011000,
	14'b10001100011001,
	14'b10001100011010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100101011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100000100,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100010101,
	14'b10010100010110,
	14'b10010100010111,
	14'b10010100011000,
	14'b10010100011001,
	14'b10010100011010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100101011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010100111011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011100010,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100010101,
	14'b10011100010110,
	14'b10011100010111,
	14'b10011100011000,
	14'b10011100011001,
	14'b10011100011010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100101011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011100111011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101001011,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10100011100001,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000: edge_mask_reg_p6[697] <= 1'b1;
 		default: edge_mask_reg_p6[697] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000000,
	14'b1101101010000,
	14'b1101101100000,
	14'b1110101000000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000: edge_mask_reg_p6[698] <= 1'b1;
 		default: edge_mask_reg_p6[698] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1111100110000,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b10000100100000,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101110000: edge_mask_reg_p6[699] <= 1'b1;
 		default: edge_mask_reg_p6[699] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110000,
	14'b10011101110001,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000: edge_mask_reg_p6[700] <= 1'b1;
 		default: edge_mask_reg_p6[700] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1111100110010,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110001,
	14'b10000101110010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110001,
	14'b10001101110010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110001,
	14'b10010101110010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110001,
	14'b10011101110010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000: edge_mask_reg_p6[701] <= 1'b1;
 		default: edge_mask_reg_p6[701] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1111100110011,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110010,
	14'b10000101110011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110010,
	14'b10001101110011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110010,
	14'b10010101110011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110010,
	14'b10011101110011,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10100101010001: edge_mask_reg_p6[702] <= 1'b1;
 		default: edge_mask_reg_p6[702] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000011,
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1111100110100,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110011,
	14'b10000101110100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110011,
	14'b10001101110100,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110011,
	14'b10010101110100,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101110011,
	14'b10011101110100,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001: edge_mask_reg_p6[703] <= 1'b1;
 		default: edge_mask_reg_p6[703] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000100,
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1110101000100,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1111100110101,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110100,
	14'b10000101110101,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110100,
	14'b10001101110101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110100,
	14'b10010101110101,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101110100,
	14'b10011101110101,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10100101010001,
	14'b10100101010010,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[704] <= 1'b1;
 		default: edge_mask_reg_p6[704] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000101,
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1110101000101,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1111100110110,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b10000011110000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110101,
	14'b10000101110110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110101,
	14'b10001101110110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110101,
	14'b10010101110110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101110101,
	14'b10011101110110,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100100100,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10101011100000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[705] <= 1'b1;
 		default: edge_mask_reg_p6[705] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000110,
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1110101000110,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100110111,
	14'b1111100111000,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110110,
	14'b10000101110111,
	14'b10001011100000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101110110,
	14'b10011101110111,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[706] <= 1'b1;
 		default: edge_mask_reg_p6[706] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101000111,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110101000111,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100111000,
	14'b1111100111001,
	14'b1111101000111,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101010000,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101110111,
	14'b10011101111000,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100011110010,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001: edge_mask_reg_p6[707] <= 1'b1;
 		default: edge_mask_reg_p6[707] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101001000,
	14'b1101101001001,
	14'b1101101001010,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1110011100000,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100110000,
	14'b1110101001000,
	14'b1110101001001,
	14'b1110101001010,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1111011100000,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100111001,
	14'b1111100111010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b10000011100000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100100111,
	14'b10000100101000,
	14'b10000100101001,
	14'b10000100101010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000100111011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10001011100000,
	14'b10001011100001,
	14'b10001011100010,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100100111,
	14'b10001100101000,
	14'b10001100101001,
	14'b10001100101010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001100111011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10010011100000,
	14'b10010011100001,
	14'b10010011100010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100100111,
	14'b10010100101000,
	14'b10010100101001,
	14'b10010100101010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010100111011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10011011100000,
	14'b10011011100001,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011011110011,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100010100,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100100110,
	14'b10011100100111,
	14'b10011100101000,
	14'b10011100101001,
	14'b10011100101010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011100111011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101001011,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101011011,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101111000,
	14'b10011101111001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001: edge_mask_reg_p6[708] <= 1'b1;
 		default: edge_mask_reg_p6[708] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010000,
	14'b1101101100000,
	14'b1101101110000,
	14'b1110101010000,
	14'b1110101100000,
	14'b1110101110000,
	14'b1111101010000,
	14'b1111101100000,
	14'b1111101110000,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10010101110001,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101110000: edge_mask_reg_p6[709] <= 1'b1;
 		default: edge_mask_reg_p6[709] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b10000100110000,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110000,
	14'b10011101110001,
	14'b10100100100000,
	14'b10100100110000: edge_mask_reg_p6[710] <= 1'b1;
 		default: edge_mask_reg_p6[710] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1111101000001,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011110000000,
	14'b10011110000001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000: edge_mask_reg_p6[711] <= 1'b1;
 		default: edge_mask_reg_p6[711] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1111101000010,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000001,
	14'b10000110000010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000001,
	14'b10001110000010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000001,
	14'b10010110000010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011110000001,
	14'b10011110000010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000: edge_mask_reg_p6[712] <= 1'b1;
 		default: edge_mask_reg_p6[712] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010010,
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1111101000011,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000010,
	14'b10000110000011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000010,
	14'b10001110000011,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000010,
	14'b10010110000011,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011110000010,
	14'b10011110000011,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001: edge_mask_reg_p6[713] <= 1'b1;
 		default: edge_mask_reg_p6[713] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010011,
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1110101010011,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1111101000100,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000011,
	14'b10000110000100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000011,
	14'b10001110000100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000011,
	14'b10010110000100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011110000011,
	14'b10011110000100,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10101011110000,
	14'b10101100000000: edge_mask_reg_p6[714] <= 1'b1;
 		default: edge_mask_reg_p6[714] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010100,
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1110101010100,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1111101000101,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000100,
	14'b10000110000101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000100,
	14'b10001110000101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000100,
	14'b10010110000101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011110000100,
	14'b10011110000101,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10100101010001,
	14'b10100101010010,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[715] <= 1'b1;
 		default: edge_mask_reg_p6[715] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010101,
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1110101010101,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1111101000110,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100100100,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000101,
	14'b10000110000110,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000101,
	14'b10001110000110,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000101,
	14'b10010110000110,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011110000101,
	14'b10011110000110,
	14'b10100011100000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100100011,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10100101010010,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[716] <= 1'b1;
 		default: edge_mask_reg_p6[716] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010110,
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1110101010110,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111101000111,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000110,
	14'b10000110000111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000110,
	14'b10001110000111,
	14'b10010011100000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010000,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000110,
	14'b10010110000111,
	14'b10011011100000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101010000,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011110000110,
	14'b10011110000111,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10101100010000,
	14'b10101100010001,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000: edge_mask_reg_p6[717] <= 1'b1;
 		default: edge_mask_reg_p6[717] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101010111,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110101010111,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100110000,
	14'b1111101001000,
	14'b1111101001001,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000111,
	14'b10000110001000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100100110,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000111,
	14'b10001110001000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000111,
	14'b10010110001000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100100,
	14'b10011100100101,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011110000111,
	14'b10011110001000,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[718] <= 1'b1;
 		default: edge_mask_reg_p6[718] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101011000,
	14'b1101101011001,
	14'b1101101011010,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100110000,
	14'b1110101000000,
	14'b1110101011000,
	14'b1110101011001,
	14'b1110101011010,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111011110010,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101001001,
	14'b1111101001010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101011000,
	14'b1111101011001,
	14'b1111101011010,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000011110011,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100100101,
	14'b10000100100110,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000100111000,
	14'b10000100111001,
	14'b10000100111010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101001011,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110001000,
	14'b10000110001001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001011110011,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000011,
	14'b10001100000100,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100100101,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001100110111,
	14'b10001100111000,
	14'b10001100111001,
	14'b10001100111010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101001011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010011110011,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100100101,
	14'b10010100100110,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010100111000,
	14'b10010100111001,
	14'b10010100111010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101001011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10011011110001,
	14'b10011011110010,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100100110,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011100110111,
	14'b10011100111000,
	14'b10011100111001,
	14'b10011100111010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101001011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101011011,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101101011,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011101111010,
	14'b10011110001000,
	14'b10011110001001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100100010,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010: edge_mask_reg_p6[719] <= 1'b1;
 		default: edge_mask_reg_p6[719] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100000,
	14'b1101101110000,
	14'b1101110000000,
	14'b1110101100000,
	14'b1110101110000,
	14'b1110110000000,
	14'b1111101100000,
	14'b1111101110000,
	14'b1111110000000,
	14'b10000101000000,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10010101000000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10010110000001,
	14'b10011101000000,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011110000000: edge_mask_reg_p6[720] <= 1'b1;
 		default: edge_mask_reg_p6[720] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110010000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011110000000,
	14'b10011110000001,
	14'b10100100110000,
	14'b10100101000000: edge_mask_reg_p6[721] <= 1'b1;
 		default: edge_mask_reg_p6[721] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10001110010001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110010000,
	14'b10010110010001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110010000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000: edge_mask_reg_p6[722] <= 1'b1;
 		default: edge_mask_reg_p6[722] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100001,
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1111101010010,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010001,
	14'b10000110010010,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010001,
	14'b10001110010010,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110010001,
	14'b10010110010010,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110010001,
	14'b10011110010010,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101100000: edge_mask_reg_p6[723] <= 1'b1;
 		default: edge_mask_reg_p6[723] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100010,
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1110101100010,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1111101010011,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b10000100110010,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010010,
	14'b10000110010011,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010010,
	14'b10001110010011,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110010010,
	14'b10010110010011,
	14'b10011100000000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110010010,
	14'b10011110010011,
	14'b10100100000000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10100101100000,
	14'b10100101100001: edge_mask_reg_p6[724] <= 1'b1;
 		default: edge_mask_reg_p6[724] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100011,
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1110101100011,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1111101010100,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b10000100110011,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010011,
	14'b10000110010100,
	14'b10001100000000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010011,
	14'b10001110010100,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110010011,
	14'b10010110010100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110010011,
	14'b10011110010100,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10100101100000,
	14'b10100101100001,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[725] <= 1'b1;
 		default: edge_mask_reg_p6[725] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100100,
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1110101100100,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1111101010101,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100110011,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010100,
	14'b10000110010101,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010100,
	14'b10001110010101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110010100,
	14'b10010110010101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110010100,
	14'b10011110010101,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100100110011,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101000011,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10100101100001,
	14'b10100101100010,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000: edge_mask_reg_p6[726] <= 1'b1;
 		default: edge_mask_reg_p6[726] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100101,
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1110101100101,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111101010110,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010101,
	14'b10000110010110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010101,
	14'b10001110010110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110010101,
	14'b10010110010110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110010101,
	14'b10011110010110,
	14'b10100011110000,
	14'b10100011110001,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100100110010,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10101011110000,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[727] <= 1'b1;
 		default: edge_mask_reg_p6[727] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101100110,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110101100110,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111101010111,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010110,
	14'b10000110010111,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010110,
	14'b10001110010111,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110010110,
	14'b10010110010111,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110010110,
	14'b10011110010111,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100000010,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100100001,
	14'b10101100110000,
	14'b10101100110001: edge_mask_reg_p6[728] <= 1'b1;
 		default: edge_mask_reg_p6[728] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101011110000,
	14'b1101100000000,
	14'b1101101100111,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110101100111,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111101000000,
	14'b1111101010000,
	14'b1111101011000,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010111,
	14'b10000110011000,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001100110110,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010111,
	14'b10001110011000,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010011110010,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100000,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110010111,
	14'b10010110011000,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100000011,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011100110100,
	14'b10011100110101,
	14'b10011100110110,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011101111010,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110001001,
	14'b10011110010111,
	14'b10011110011000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[729] <= 1'b1;
 		default: edge_mask_reg_p6[729] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100100000000,
	14'b1101011110000,
	14'b1101011110001,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101101101000,
	14'b1101101101001,
	14'b1101101101010,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1110011110000,
	14'b1110011110001,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101101000,
	14'b1110101101001,
	14'b1110101101010,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1111011110000,
	14'b1111011110001,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101011001,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101101010,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b10000011110000,
	14'b10000011110001,
	14'b10000011110010,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000100110110,
	14'b10000100110111,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101001000,
	14'b10000101001001,
	14'b10000101001010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101011011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110011000,
	14'b10000110011001,
	14'b10001011110000,
	14'b10001011110001,
	14'b10001011110010,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101001000,
	14'b10001101001001,
	14'b10001101001010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101011011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110011000,
	14'b10001110011001,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100000011,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100010100,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100100100,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010100110101,
	14'b10010100110110,
	14'b10010100110111,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101001000,
	14'b10010101001001,
	14'b10010101001010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101011011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010101111011,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110011000,
	14'b10010110011001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000110,
	14'b10011101000111,
	14'b10011101001000,
	14'b10011101001001,
	14'b10011101001010,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101011011,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101101011,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011101111010,
	14'b10011101111011,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110001001,
	14'b10011110001010,
	14'b10011110011000,
	14'b10011110011001: edge_mask_reg_p6[730] <= 1'b1;
 		default: edge_mask_reg_p6[730] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110000,
	14'b1101110000000,
	14'b1101110010000,
	14'b1110101110000,
	14'b1110110000000,
	14'b1110110010000,
	14'b1111101110000,
	14'b1111110000000,
	14'b1111110010000,
	14'b10000101010000,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110010000,
	14'b10000110010001,
	14'b10001101010000,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110010000,
	14'b10001110010001,
	14'b10010101010000,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110010000,
	14'b10010110010001,
	14'b10011101010000,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110010000,
	14'b10100101010000: edge_mask_reg_p6[731] <= 1'b1;
 		default: edge_mask_reg_p6[731] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110000,
	14'b1101101110001,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110010000,
	14'b1101110010001,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110010000,
	14'b1110110010001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110010000,
	14'b1111110010001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10001101000000,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110100000,
	14'b10010101000000,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110010000,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110100000,
	14'b10011101000000,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110010000,
	14'b10011110010001,
	14'b10100101000000,
	14'b10100101010000: edge_mask_reg_p6[732] <= 1'b1;
 		default: edge_mask_reg_p6[732] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110000,
	14'b1101101110001,
	14'b1101101110010,
	14'b1101110000000,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110010000,
	14'b1101110010001,
	14'b1101110010010,
	14'b1110101110000,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110110000000,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110010000,
	14'b1110110010001,
	14'b1110110010010,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111110000000,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110010000,
	14'b1111110010001,
	14'b1111110010010,
	14'b10000101000001,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110100000,
	14'b10000110100001,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110100000,
	14'b10001110100001,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110010000,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110100000,
	14'b10010110100001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110010000,
	14'b10011110010001,
	14'b10011110010010,
	14'b10011110100000,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101100000: edge_mask_reg_p6[733] <= 1'b1;
 		default: edge_mask_reg_p6[733] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110001,
	14'b1101101110010,
	14'b1101101110011,
	14'b1101110000001,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110010001,
	14'b1101110010010,
	14'b1101110010011,
	14'b1110101110001,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110110000001,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110010001,
	14'b1110110010010,
	14'b1110110010011,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111110000001,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110010001,
	14'b1111110010010,
	14'b1111110010011,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110010000,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110100001,
	14'b10000110100010,
	14'b10001100110000,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110010000,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110100001,
	14'b10001110100010,
	14'b10010100110000,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110010000,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110100001,
	14'b10010110100010,
	14'b10011100010000,
	14'b10011100110000,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110010000,
	14'b10011110010001,
	14'b10011110010010,
	14'b10011110010011,
	14'b10011110100001,
	14'b10100100010000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101100000,
	14'b10100101100001,
	14'b10100101110000: edge_mask_reg_p6[734] <= 1'b1;
 		default: edge_mask_reg_p6[734] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110010,
	14'b1101101110011,
	14'b1101101110100,
	14'b1101110000010,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110010010,
	14'b1101110010011,
	14'b1101110010100,
	14'b1110101110010,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110110000010,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110010010,
	14'b1110110010011,
	14'b1110110010100,
	14'b1111101110010,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111110000010,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110010010,
	14'b1111110010011,
	14'b1111110010100,
	14'b10000101000010,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000110000000,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110010001,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110100010,
	14'b10000110100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001110000000,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110010001,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110100010,
	14'b10001110100011,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010110000000,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110010001,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110100010,
	14'b10010110100011,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011110000000,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110010001,
	14'b10011110010010,
	14'b10011110010011,
	14'b10011110010100,
	14'b10011110100010,
	14'b10011110100011,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10100101100000,
	14'b10100101100001,
	14'b10100101110000,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[735] <= 1'b1;
 		default: edge_mask_reg_p6[735] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110011,
	14'b1101101110100,
	14'b1101101110101,
	14'b1101110000011,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110010011,
	14'b1101110010100,
	14'b1101110010101,
	14'b1110101110011,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110110000011,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110010011,
	14'b1110110010100,
	14'b1110110010101,
	14'b1111101100100,
	14'b1111101110011,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111110000011,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110010011,
	14'b1111110010100,
	14'b1111110010101,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000110000001,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110010010,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110100011,
	14'b10000110100100,
	14'b10001100000000,
	14'b10001100010000,
	14'b10001100100000,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101110000,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001110000001,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110010010,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110100011,
	14'b10001110100100,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101110000,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010110000001,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110010010,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110100011,
	14'b10010110100100,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101110000,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011110000001,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110010010,
	14'b10011110010011,
	14'b10011110010100,
	14'b10011110010101,
	14'b10011110100011,
	14'b10011110100100,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10100101100000,
	14'b10100101100001,
	14'b10100101100010,
	14'b10101100000000,
	14'b10101100010000: edge_mask_reg_p6[736] <= 1'b1;
 		default: edge_mask_reg_p6[736] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110100,
	14'b1101101110101,
	14'b1101101110110,
	14'b1101110000100,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110010100,
	14'b1101110010101,
	14'b1101110010110,
	14'b1110101110100,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110110000100,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110010100,
	14'b1110110010101,
	14'b1110110010110,
	14'b1111100000000,
	14'b1111101100101,
	14'b1111101110100,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111110000100,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110010100,
	14'b1111110010101,
	14'b1111110010110,
	14'b10000100000000,
	14'b10000100010000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101110001,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000110000010,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110010011,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110100100,
	14'b10000110100101,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101110001,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001110000010,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110010011,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110100100,
	14'b10001110100101,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101110001,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010110000010,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110010011,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110100100,
	14'b10010110100101,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101100000,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101110001,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011110000010,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110010011,
	14'b10011110010100,
	14'b10011110010101,
	14'b10011110010110,
	14'b10011110100100,
	14'b10011110100101,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101000010,
	14'b10100101010000,
	14'b10100101010001,
	14'b10100101010010,
	14'b10101100000000,
	14'b10101100010000,
	14'b10101100100000,
	14'b10101100110000: edge_mask_reg_p6[737] <= 1'b1;
 		default: edge_mask_reg_p6[737] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110101,
	14'b1101101110110,
	14'b1101101110111,
	14'b1101110000101,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110010101,
	14'b1101110010110,
	14'b1101110010111,
	14'b1110100000000,
	14'b1110101110101,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110110000101,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110010101,
	14'b1110110010110,
	14'b1110110010111,
	14'b1111100000000,
	14'b1111100010000,
	14'b1111101100110,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110010101,
	14'b1111110010110,
	14'b1111110010111,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100110000,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101110010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000110000011,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110010100,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110100101,
	14'b10000110100110,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101110010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001110000011,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110010100,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110100101,
	14'b10001110100110,
	14'b10010011110000,
	14'b10010011110001,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101110010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010110000011,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110010100,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110100101,
	14'b10010110100110,
	14'b10011011110000,
	14'b10011011110001,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101100001,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101110010,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011110000011,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110010100,
	14'b10011110010101,
	14'b10011110010110,
	14'b10011110010111,
	14'b10011110100101,
	14'b10011110100110,
	14'b10100011110000,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001,
	14'b10100101010000,
	14'b10101100100000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[738] <= 1'b1;
 		default: edge_mask_reg_p6[738] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101101110110,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101110000110,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110010110,
	14'b1101110010111,
	14'b1101110011000,
	14'b1110100000000,
	14'b1110100010000,
	14'b1110101110110,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110110000110,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110010110,
	14'b1110110010111,
	14'b1110110011000,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111101100111,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110010110,
	14'b1111110010111,
	14'b1111110011000,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110010101,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110100110,
	14'b10000110100111,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110010101,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110100110,
	14'b10001110100111,
	14'b10010011110000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110010101,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110100110,
	14'b10010110100111,
	14'b10011011110000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011100110011,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010010,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101100000,
	14'b10011101100010,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101110011,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110001001,
	14'b10011110010101,
	14'b10011110010110,
	14'b10011110010111,
	14'b10011110011000,
	14'b10011110100110,
	14'b10011110100111,
	14'b10100100000000,
	14'b10100100000001,
	14'b10100100010000,
	14'b10100100010001,
	14'b10100100010010,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10101100110000,
	14'b10101101000000: edge_mask_reg_p6[739] <= 1'b1;
 		default: edge_mask_reg_p6[739] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1101100000000,
	14'b1101100010000,
	14'b1101101110111,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101110000111,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110010111,
	14'b1101110011000,
	14'b1101110011001,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110101110111,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110110000111,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110010111,
	14'b1110110011000,
	14'b1110110011001,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101100000,
	14'b1111101101000,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110010111,
	14'b1111110011000,
	14'b1111110011001,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101110011,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000110000100,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110010110,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110100111,
	14'b10000110101000,
	14'b10001011110000,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101110011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001110000100,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110100111,
	14'b10001110101000,
	14'b10010100000000,
	14'b10010100000001,
	14'b10010100000010,
	14'b10010100010000,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010100110100,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000100,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010011,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100010,
	14'b10010101100011,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101110011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010110000100,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110010110,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110011001,
	14'b10010110100111,
	14'b10010110101000,
	14'b10011100000000,
	14'b10011100000001,
	14'b10011100000010,
	14'b10011100010000,
	14'b10011100010001,
	14'b10011100010010,
	14'b10011100010011,
	14'b10011100100000,
	14'b10011100100001,
	14'b10011100100010,
	14'b10011100100011,
	14'b10011100110000,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000000,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101000011,
	14'b10011101000100,
	14'b10011101000101,
	14'b10011101000110,
	14'b10011101010000,
	14'b10011101010001,
	14'b10011101010011,
	14'b10011101010100,
	14'b10011101010101,
	14'b10011101010110,
	14'b10011101010111,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101100000,
	14'b10011101100011,
	14'b10011101100100,
	14'b10011101100101,
	14'b10011101100110,
	14'b10011101100111,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101110100,
	14'b10011101110101,
	14'b10011101110110,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011101111010,
	14'b10011110000100,
	14'b10011110000101,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110001001,
	14'b10011110001010,
	14'b10011110010110,
	14'b10011110010111,
	14'b10011110011000,
	14'b10011110011001,
	14'b10011110100111,
	14'b10011110101000,
	14'b10100100100000,
	14'b10100100100001,
	14'b10100100110000,
	14'b10100100110001,
	14'b10100101000000,
	14'b10100101000001: edge_mask_reg_p6[740] <= 1'b1;
 		default: edge_mask_reg_p6[740] <= 1'b0;
 	endcase

    case({z,y,x})
	14'b1100011110000,
	14'b1100100000000,
	14'b1100100000001,
	14'b1100100010000,
	14'b1100100010001,
	14'b1101011110000,
	14'b1101100000000,
	14'b1101100000001,
	14'b1101100000010,
	14'b1101100010000,
	14'b1101100010001,
	14'b1101100010010,
	14'b1101100010011,
	14'b1101100100000,
	14'b1101100100001,
	14'b1101100100010,
	14'b1101100100011,
	14'b1101100110000,
	14'b1101100110001,
	14'b1101100110010,
	14'b1101100110011,
	14'b1101101000000,
	14'b1101101000001,
	14'b1101101000010,
	14'b1101101000011,
	14'b1101101010000,
	14'b1101101010001,
	14'b1101101010010,
	14'b1101101100000,
	14'b1101101100001,
	14'b1101101111000,
	14'b1101101111001,
	14'b1101101111010,
	14'b1101110001000,
	14'b1101110001001,
	14'b1101110001010,
	14'b1101110011000,
	14'b1101110011001,
	14'b1101110011010,
	14'b1110011110000,
	14'b1110100000000,
	14'b1110100000001,
	14'b1110100000010,
	14'b1110100000011,
	14'b1110100010000,
	14'b1110100010001,
	14'b1110100010010,
	14'b1110100010011,
	14'b1110100010100,
	14'b1110100100000,
	14'b1110100100001,
	14'b1110100100010,
	14'b1110100100011,
	14'b1110100100100,
	14'b1110100110000,
	14'b1110100110001,
	14'b1110100110010,
	14'b1110100110011,
	14'b1110100110100,
	14'b1110101000000,
	14'b1110101000001,
	14'b1110101000010,
	14'b1110101000011,
	14'b1110101000100,
	14'b1110101010000,
	14'b1110101010001,
	14'b1110101010010,
	14'b1110101010011,
	14'b1110101100000,
	14'b1110101100001,
	14'b1110101100010,
	14'b1110101110000,
	14'b1110101111000,
	14'b1110101111001,
	14'b1110101111010,
	14'b1110110001000,
	14'b1110110001001,
	14'b1110110001010,
	14'b1110110011000,
	14'b1110110011001,
	14'b1110110011010,
	14'b1111011110000,
	14'b1111100000000,
	14'b1111100000001,
	14'b1111100000010,
	14'b1111100000011,
	14'b1111100010000,
	14'b1111100010001,
	14'b1111100010010,
	14'b1111100010011,
	14'b1111100010100,
	14'b1111100100000,
	14'b1111100100001,
	14'b1111100100010,
	14'b1111100100011,
	14'b1111100100100,
	14'b1111100110000,
	14'b1111100110001,
	14'b1111100110010,
	14'b1111100110011,
	14'b1111100110100,
	14'b1111100110101,
	14'b1111101000000,
	14'b1111101000001,
	14'b1111101000010,
	14'b1111101000011,
	14'b1111101000100,
	14'b1111101000101,
	14'b1111101000110,
	14'b1111101000111,
	14'b1111101010000,
	14'b1111101010001,
	14'b1111101010010,
	14'b1111101010011,
	14'b1111101010100,
	14'b1111101010101,
	14'b1111101010110,
	14'b1111101010111,
	14'b1111101011000,
	14'b1111101100000,
	14'b1111101100001,
	14'b1111101100010,
	14'b1111101100011,
	14'b1111101100100,
	14'b1111101100101,
	14'b1111101100110,
	14'b1111101100111,
	14'b1111101101000,
	14'b1111101101001,
	14'b1111101110000,
	14'b1111101110001,
	14'b1111101110010,
	14'b1111101110101,
	14'b1111101110110,
	14'b1111101110111,
	14'b1111101111000,
	14'b1111101111001,
	14'b1111101111010,
	14'b1111110000101,
	14'b1111110000110,
	14'b1111110000111,
	14'b1111110001000,
	14'b1111110001001,
	14'b1111110001010,
	14'b1111110011000,
	14'b1111110011001,
	14'b1111110011010,
	14'b10000011110000,
	14'b10000100000000,
	14'b10000100000001,
	14'b10000100000010,
	14'b10000100000011,
	14'b10000100010000,
	14'b10000100010001,
	14'b10000100010010,
	14'b10000100010011,
	14'b10000100010100,
	14'b10000100100000,
	14'b10000100100001,
	14'b10000100100010,
	14'b10000100100011,
	14'b10000100100100,
	14'b10000100110000,
	14'b10000100110001,
	14'b10000100110010,
	14'b10000100110011,
	14'b10000100110100,
	14'b10000100110101,
	14'b10000101000000,
	14'b10000101000001,
	14'b10000101000010,
	14'b10000101000011,
	14'b10000101000100,
	14'b10000101000101,
	14'b10000101000110,
	14'b10000101000111,
	14'b10000101010000,
	14'b10000101010001,
	14'b10000101010010,
	14'b10000101010011,
	14'b10000101010100,
	14'b10000101010101,
	14'b10000101010110,
	14'b10000101010111,
	14'b10000101011000,
	14'b10000101011001,
	14'b10000101011010,
	14'b10000101100000,
	14'b10000101100001,
	14'b10000101100010,
	14'b10000101100011,
	14'b10000101100100,
	14'b10000101100101,
	14'b10000101100110,
	14'b10000101100111,
	14'b10000101101000,
	14'b10000101101001,
	14'b10000101101010,
	14'b10000101101011,
	14'b10000101110000,
	14'b10000101110001,
	14'b10000101110100,
	14'b10000101110101,
	14'b10000101110110,
	14'b10000101110111,
	14'b10000101111000,
	14'b10000101111001,
	14'b10000101111010,
	14'b10000101111011,
	14'b10000110000101,
	14'b10000110000110,
	14'b10000110000111,
	14'b10000110001000,
	14'b10000110001001,
	14'b10000110001010,
	14'b10000110001011,
	14'b10000110010111,
	14'b10000110011000,
	14'b10000110011001,
	14'b10000110011010,
	14'b10000110101000,
	14'b10000110101001,
	14'b10001100000000,
	14'b10001100000001,
	14'b10001100000010,
	14'b10001100000011,
	14'b10001100010000,
	14'b10001100010001,
	14'b10001100010010,
	14'b10001100010011,
	14'b10001100010100,
	14'b10001100100000,
	14'b10001100100001,
	14'b10001100100010,
	14'b10001100100011,
	14'b10001100100100,
	14'b10001100110000,
	14'b10001100110001,
	14'b10001100110010,
	14'b10001100110011,
	14'b10001100110100,
	14'b10001100110101,
	14'b10001101000000,
	14'b10001101000001,
	14'b10001101000010,
	14'b10001101000011,
	14'b10001101000100,
	14'b10001101000101,
	14'b10001101000110,
	14'b10001101000111,
	14'b10001101010000,
	14'b10001101010001,
	14'b10001101010010,
	14'b10001101010011,
	14'b10001101010100,
	14'b10001101010101,
	14'b10001101010110,
	14'b10001101010111,
	14'b10001101011000,
	14'b10001101011001,
	14'b10001101011010,
	14'b10001101100000,
	14'b10001101100001,
	14'b10001101100010,
	14'b10001101100011,
	14'b10001101100100,
	14'b10001101100101,
	14'b10001101100110,
	14'b10001101100111,
	14'b10001101101000,
	14'b10001101101001,
	14'b10001101101010,
	14'b10001101101011,
	14'b10001101110100,
	14'b10001101110101,
	14'b10001101110110,
	14'b10001101110111,
	14'b10001101111000,
	14'b10001101111001,
	14'b10001101111010,
	14'b10001101111011,
	14'b10001110000101,
	14'b10001110000110,
	14'b10001110000111,
	14'b10001110001000,
	14'b10001110001001,
	14'b10001110001010,
	14'b10001110001011,
	14'b10001110010110,
	14'b10001110010111,
	14'b10001110011000,
	14'b10001110011001,
	14'b10001110011010,
	14'b10001110101000,
	14'b10001110101001,
	14'b10010100000010,
	14'b10010100010001,
	14'b10010100010010,
	14'b10010100010011,
	14'b10010100100000,
	14'b10010100100001,
	14'b10010100100010,
	14'b10010100100011,
	14'b10010100110000,
	14'b10010100110001,
	14'b10010100110010,
	14'b10010100110011,
	14'b10010101000000,
	14'b10010101000001,
	14'b10010101000010,
	14'b10010101000011,
	14'b10010101000101,
	14'b10010101000110,
	14'b10010101000111,
	14'b10010101010000,
	14'b10010101010001,
	14'b10010101010010,
	14'b10010101010100,
	14'b10010101010101,
	14'b10010101010110,
	14'b10010101010111,
	14'b10010101011000,
	14'b10010101011001,
	14'b10010101011010,
	14'b10010101100000,
	14'b10010101100001,
	14'b10010101100100,
	14'b10010101100101,
	14'b10010101100110,
	14'b10010101100111,
	14'b10010101101000,
	14'b10010101101001,
	14'b10010101101010,
	14'b10010101101011,
	14'b10010101110100,
	14'b10010101110101,
	14'b10010101110110,
	14'b10010101110111,
	14'b10010101111000,
	14'b10010101111001,
	14'b10010101111010,
	14'b10010101111011,
	14'b10010110000101,
	14'b10010110000110,
	14'b10010110000111,
	14'b10010110001000,
	14'b10010110001001,
	14'b10010110001010,
	14'b10010110001011,
	14'b10010110010111,
	14'b10010110011000,
	14'b10010110011001,
	14'b10010110011010,
	14'b10010110101000,
	14'b10010110101001,
	14'b10011100110001,
	14'b10011100110010,
	14'b10011101000001,
	14'b10011101000010,
	14'b10011101011000,
	14'b10011101011001,
	14'b10011101011010,
	14'b10011101101000,
	14'b10011101101001,
	14'b10011101101010,
	14'b10011101101011,
	14'b10011101110111,
	14'b10011101111000,
	14'b10011101111001,
	14'b10011101111010,
	14'b10011101111011,
	14'b10011110000110,
	14'b10011110000111,
	14'b10011110001000,
	14'b10011110001001,
	14'b10011110001010,
	14'b10011110001011,
	14'b10011110010111,
	14'b10011110011000,
	14'b10011110011001,
	14'b10011110011010,
	14'b10011110101000,
	14'b10011110101001,
	14'b10100101111001,
	14'b10100101111010,
	14'b10100110001001: edge_mask_reg_p6[741] <= 1'b1;
 		default: edge_mask_reg_p6[741] <= 1'b0;
 	endcase

end
endmodule

