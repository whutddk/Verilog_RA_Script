
`timescale 1 ns / 1 ns

////////////////////////////////////////////////////////////////////////////////
// Company: Wuhan university of technology 
// Engineer: Ruige LEE
//
// Create Date: 20181202
// Design Name: pkb-2019
// Module Name: flatten
// Target Device: <zynq7000-z020>
// Tool versions: <2018.02>
// Description:
//    
// Dependencies:
//    
// Revision:
//    0.1.0
// Additional Comments:
//    
////////////////////////////////////////////////////////////////////////////////
			

module graph
(

)


//state Ram:0-1024
always @(posedge CLK or !RST_n) begin
	if (!RST_n) begin
		// reset
		
	end
	else if () begin
		
	end
end


//state lever 0-10
always @(posedge CLK or !RST_n) begin
	if (!RST_n) begin
		// reset
		
	end
	else if () begin
		
	end
end



//state INIT FORWARD BACKWARD 
always @(negedge CLK or !RST_n) begin
	if (!RST_n) begin
		// reset
		
	end
	else if ( state == INIT ) begin
		maxLever <= 4'D10;
		ActivePose <= (65'b1 << startPoint);
		edgeMask_reg[1033:0] <= edgeMask[1033:0];

		edgeActive[0] <= 1034'b0;
		edgeActive[1] <= 1034'b0;
		edgeActive[2] <= 1034'b0;
		edgeActive[3] <= 1034'b0;
		edgeActive[4] <= 1034'b0;
		edgeActive[5] <= 1034'b0;
		edgeActive[6] <= 1034'b0;
		edgeActive[7] <= 1034'b0;
		edgeActive[8] <= 1034'b0;
		edgeActive[9] <= 1034'b0;


		// RAM_address <= 10'd0;

	end

	else if (state == FORWARD) begin
		


		if( (ActivePose >> endpoint) & 1'B1 == 1 ) begin
			state <= BACKWARD;
			edgeMask_reg <= edgeMask_reg 
							| edgeActive[0] | edgeActive[1] | edgeActive[2] | edgeActive[3]
							| edgeActive[4] | edgeActive[5] | edgeActive[6] | edgeActive[7]
							| edgeActive[8] | edgeActive[9] ;
			maxLever <= poseLeverCnt
			ActivePose <= (65'b1 << ENDPoint);
		end

		else begin
			state <= FORWARD;
		end

	end

	else if ( state == c )begin
		
	end

	else begin//idle


	end


end

endmodule

