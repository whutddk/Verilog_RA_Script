/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 5
second: 57
********************************************/

module prm_LUTX1_Sp_4_4_4_chk512p3(
	input [3:0] x,
	input [3:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p3
);

	reg [511:0] edge_mask_reg_512p3;
	assign edge_mask_512p3= edge_mask_reg_512p3;

always @( *) begin
    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101101110100,
12'b101110000100,
12'b101110010100: edge_mask_reg_512p3[0] <= 1'b1;
 		default: edge_mask_reg_512p3[0] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b101001000100,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101101000100,
12'b101101010100,
12'b101101100100: edge_mask_reg_512p3[1] <= 1'b1;
 		default: edge_mask_reg_512p3[1] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101101000100,
12'b101101010100,
12'b101101100100: edge_mask_reg_512p3[2] <= 1'b1;
 		default: edge_mask_reg_512p3[2] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101101000100,
12'b101101010100,
12'b101101100100: edge_mask_reg_512p3[3] <= 1'b1;
 		default: edge_mask_reg_512p3[3] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100101010,
12'b10100110110,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b100000110101,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101101000100,
12'b101101000101,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b110001000100: edge_mask_reg_512p3[4] <= 1'b1;
 		default: edge_mask_reg_512p3[4] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100101010,
12'b10100110110,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000110101,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101101000100,
12'b101101000101,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b110001000100: edge_mask_reg_512p3[5] <= 1'b1;
 		default: edge_mask_reg_512p3[5] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101001110100: edge_mask_reg_512p3[6] <= 1'b1;
 		default: edge_mask_reg_512p3[6] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010010011: edge_mask_reg_512p3[7] <= 1'b1;
 		default: edge_mask_reg_512p3[7] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[8] <= 1'b1;
 		default: edge_mask_reg_512p3[8] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[9] <= 1'b1;
 		default: edge_mask_reg_512p3[9] <= 1'b0;
 	endcase

    case({x,y,z})
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011010111,
12'b1011011000,
12'b1011011001,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10011001000,
12'b10011001001,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10111001000,
12'b10111001001,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11111011000,
12'b11111011001,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011110110,
12'b100011110111,
12'b100111010110,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110101,
12'b100111110110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011110101,
12'b101011110110,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111110100,
12'b101111110101,
12'b101111110110,
12'b110011100100,
12'b110011100101,
12'b110011100110,
12'b110011110100,
12'b110011110101,
12'b110011110110,
12'b110111100100,
12'b110111100101,
12'b110111110100,
12'b110111110101,
12'b111011100100,
12'b111011110100: edge_mask_reg_512p3[10] <= 1'b1;
 		default: edge_mask_reg_512p3[10] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011010111,
12'b1011011000,
12'b1011011001,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11111001000,
12'b11111001001,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011110110,
12'b100011110111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110101,
12'b100111110110,
12'b100111110111,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011110101,
12'b101011110110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111110100,
12'b101111110101,
12'b101111110110,
12'b110011010100,
12'b110011010101,
12'b110011010110,
12'b110011100100,
12'b110011100101,
12'b110011100110,
12'b110011110100,
12'b110011110101,
12'b110011110110,
12'b110111010100,
12'b110111100100,
12'b110111110100: edge_mask_reg_512p3[11] <= 1'b1;
 		default: edge_mask_reg_512p3[11] <= 1'b0;
 	endcase

    case({x,y,z})
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011010111,
12'b1011011000,
12'b1011011001,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10011001000,
12'b10011001001,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10111001000,
12'b10111001001,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11111011000,
12'b11111011001,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011110110,
12'b100011110111,
12'b100111010110,
12'b100111100101,
12'b100111100110,
12'b100111110101,
12'b100111110110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011110101,
12'b101011110110,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111110100,
12'b101111110101,
12'b101111110110,
12'b110011100100,
12'b110011100101,
12'b110011100110,
12'b110011110100,
12'b110011110101,
12'b110011110110,
12'b110111100100,
12'b110111110100: edge_mask_reg_512p3[12] <= 1'b1;
 		default: edge_mask_reg_512p3[12] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110101,
12'b1110110,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000101,
12'b10000110,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10001001001,
12'b10001001010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10101001001,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001010100,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001001,
12'b11110001010,
12'b100001100011,
12'b100001110011,
12'b100001110100,
12'b100010000011: edge_mask_reg_512p3[13] <= 1'b1;
 		default: edge_mask_reg_512p3[13] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1000110111,
12'b1000111000,
12'b1000111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010101,
12'b101001010110,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101101000101,
12'b101101000110,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110101000100,
12'b110101000101,
12'b110101000110,
12'b110101010100,
12'b110101010101,
12'b110101010110,
12'b110101100100,
12'b110101100101,
12'b110101100110,
12'b111001000100,
12'b111001000101,
12'b111001010100,
12'b111001010101,
12'b111001100100,
12'b111001100101,
12'b111101010101: edge_mask_reg_512p3[14] <= 1'b1;
 		default: edge_mask_reg_512p3[14] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001001,
12'b11001001010,
12'b11001011001,
12'b11001011010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000101,
12'b100001000110,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000101,
12'b100101000110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100100100,
12'b101100100101,
12'b101100110100,
12'b101100110101,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000110100,
12'b110000110101: edge_mask_reg_512p3[15] <= 1'b1;
 		default: edge_mask_reg_512p3[15] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101001001,
12'b11101001010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100100100,
12'b101100100101,
12'b101100110100,
12'b101100110101,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000110101: edge_mask_reg_512p3[16] <= 1'b1;
 		default: edge_mask_reg_512p3[16] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101: edge_mask_reg_512p3[17] <= 1'b1;
 		default: edge_mask_reg_512p3[17] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101001000110,
12'b101100010100,
12'b101100010101,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000100110,
12'b110000110100,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[18] <= 1'b1;
 		default: edge_mask_reg_512p3[18] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100100,
12'b101001100101,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100100,
12'b101101100101,
12'b110001000101,
12'b110001010100,
12'b110001010101: edge_mask_reg_512p3[19] <= 1'b1;
 		default: edge_mask_reg_512p3[19] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111010,
12'b11110111011,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100110001000,
12'b100110001001,
12'b100110011000,
12'b100110011001,
12'b100110011010,
12'b100110101000,
12'b100110101001,
12'b100110101010,
12'b101010001000,
12'b101010001001,
12'b101010011000,
12'b101010011001,
12'b101010101000,
12'b101010101001,
12'b101110000111,
12'b101110001000,
12'b101110001001,
12'b101110010111,
12'b101110011000,
12'b101110011001,
12'b101110101000,
12'b101110101001,
12'b110010000111,
12'b110010001000,
12'b110010001001,
12'b110010010111,
12'b110010011000,
12'b110010011001,
12'b110010101000,
12'b110010101001,
12'b110110000111,
12'b110110001000,
12'b110110001001,
12'b110110010111,
12'b110110011000,
12'b110110011001,
12'b110110100111,
12'b110110101000,
12'b110110101001,
12'b111010000111,
12'b111010001000,
12'b111010010111,
12'b111010011000,
12'b111010011001,
12'b111010100111,
12'b111010101000,
12'b111110000111,
12'b111110001000,
12'b111110010111,
12'b111110011000,
12'b111110100111: edge_mask_reg_512p3[20] <= 1'b1;
 		default: edge_mask_reg_512p3[20] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110101,
12'b101010110110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110110010100,
12'b110110010101,
12'b110110100100,
12'b110110100101: edge_mask_reg_512p3[21] <= 1'b1;
 		default: edge_mask_reg_512p3[21] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110000111,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111110010110,
12'b111110010111,
12'b111110100110: edge_mask_reg_512p3[22] <= 1'b1;
 		default: edge_mask_reg_512p3[22] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100110000111,
12'b100110001000,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110000111,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111110010110,
12'b111110010111,
12'b111110100110: edge_mask_reg_512p3[23] <= 1'b1;
 		default: edge_mask_reg_512p3[23] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101010,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111010,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101: edge_mask_reg_512p3[24] <= 1'b1;
 		default: edge_mask_reg_512p3[24] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010101: edge_mask_reg_512p3[25] <= 1'b1;
 		default: edge_mask_reg_512p3[25] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111010,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b101001010101,
12'b101001010110,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b110001010101,
12'b110001100101,
12'b110001110101: edge_mask_reg_512p3[26] <= 1'b1;
 		default: edge_mask_reg_512p3[26] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100111000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100: edge_mask_reg_512p3[27] <= 1'b1;
 		default: edge_mask_reg_512p3[27] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100: edge_mask_reg_512p3[28] <= 1'b1;
 		default: edge_mask_reg_512p3[28] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101110100100,
12'b101110110100: edge_mask_reg_512p3[29] <= 1'b1;
 		default: edge_mask_reg_512p3[29] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100111000011,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100: edge_mask_reg_512p3[30] <= 1'b1;
 		default: edge_mask_reg_512p3[30] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010010101,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010100,
12'b10111010101,
12'b10111010110,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010100,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010101,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101011000011,
12'b101011000100,
12'b101110110100: edge_mask_reg_512p3[31] <= 1'b1;
 		default: edge_mask_reg_512p3[31] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101110010100,
12'b101110100100,
12'b101110110100: edge_mask_reg_512p3[32] <= 1'b1;
 		default: edge_mask_reg_512p3[32] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101000,
12'b10011101001,
12'b10110001001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101000,
12'b11011101001,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111011000,
12'b11111011001,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010100,
12'b100011010101,
12'b100011010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010011,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010011,
12'b101011010100,
12'b101011010101,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110110100,
12'b110110110101,
12'b110111000100,
12'b110111000101: edge_mask_reg_512p3[33] <= 1'b1;
 		default: edge_mask_reg_512p3[33] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110101,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000101,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010110,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101100100,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110101,
12'b110110110,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001100100,
12'b1001100101,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001100100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010001010,
12'b100010011010: edge_mask_reg_512p3[34] <= 1'b1;
 		default: edge_mask_reg_512p3[34] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100101,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110100101,
12'b111010000101,
12'b111010000110,
12'b111010010101: edge_mask_reg_512p3[35] <= 1'b1;
 		default: edge_mask_reg_512p3[35] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010100100: edge_mask_reg_512p3[36] <= 1'b1;
 		default: edge_mask_reg_512p3[36] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010100100: edge_mask_reg_512p3[37] <= 1'b1;
 		default: edge_mask_reg_512p3[37] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010100100: edge_mask_reg_512p3[38] <= 1'b1;
 		default: edge_mask_reg_512p3[38] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010100100: edge_mask_reg_512p3[39] <= 1'b1;
 		default: edge_mask_reg_512p3[39] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001100110,
12'b11001100111,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101100101,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100110,
12'b100110100111,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110: edge_mask_reg_512p3[40] <= 1'b1;
 		default: edge_mask_reg_512p3[40] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001100110,
12'b11001100111,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100110,
12'b100110100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110: edge_mask_reg_512p3[41] <= 1'b1;
 		default: edge_mask_reg_512p3[41] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001100111,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100110,
12'b100110100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101101110101,
12'b101101110110,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110: edge_mask_reg_512p3[42] <= 1'b1;
 		default: edge_mask_reg_512p3[42] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100111,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010110,
12'b100110010111,
12'b100110100110,
12'b100110100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110: edge_mask_reg_512p3[43] <= 1'b1;
 		default: edge_mask_reg_512p3[43] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001101010,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001111010,
12'b100010000100,
12'b100010000101,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b101001100100,
12'b101001100101,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101: edge_mask_reg_512p3[44] <= 1'b1;
 		default: edge_mask_reg_512p3[44] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101010,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010101,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101: edge_mask_reg_512p3[45] <= 1'b1;
 		default: edge_mask_reg_512p3[45] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100110,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011001,
12'b11011011010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100111000011,
12'b100111000100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101011000011,
12'b101011000100: edge_mask_reg_512p3[46] <= 1'b1;
 		default: edge_mask_reg_512p3[46] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111010,
12'b10110111011,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111010,
12'b11010111011,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101101010,
12'b11101101011,
12'b11101101100,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110101010,
12'b11110101011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001111010,
12'b100001111011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010001010,
12'b100010001011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b101001110101,
12'b101010000101,
12'b101010010101: edge_mask_reg_512p3[47] <= 1'b1;
 		default: edge_mask_reg_512p3[47] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001010,
12'b100111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100101000,
12'b1100101001,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111010,
12'b1101111011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100101001,
12'b11100101010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100100110011,
12'b100100110100,
12'b100101000011,
12'b100101000100,
12'b100101010011,
12'b100101010100,
12'b101000110011,
12'b101000110100,
12'b101001000011,
12'b101001000100,
12'b101001010011,
12'b101001010100: edge_mask_reg_512p3[48] <= 1'b1;
 		default: edge_mask_reg_512p3[48] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b100111000,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b1000110110,
12'b1000110111,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b10000100101,
12'b10000100110,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11100100100,
12'b11100100101,
12'b11100101001,
12'b11100101010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b100000110011,
12'b100000110100,
12'b100001000011,
12'b100001000100,
12'b100001010011,
12'b100001010100,
12'b100100110011,
12'b100100110100,
12'b100101000011,
12'b100101000100,
12'b100101010011,
12'b100101010100,
12'b101000110011,
12'b101001000011: edge_mask_reg_512p3[49] <= 1'b1;
 		default: edge_mask_reg_512p3[49] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001010,
12'b100111000,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000110111,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111001,
12'b1101111010,
12'b10000100101,
12'b10000100110,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111001,
12'b10001111010,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100100100,
12'b11100100101,
12'b11100101001,
12'b11100101010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100100,
12'b100001100101,
12'b100100110011,
12'b100100110100,
12'b100101000011,
12'b100101000100,
12'b100101010011,
12'b100101010100,
12'b101000110011,
12'b101000110100,
12'b101001000011,
12'b101001000100,
12'b101001010011,
12'b101001010100: edge_mask_reg_512p3[50] <= 1'b1;
 		default: edge_mask_reg_512p3[50] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111000,
12'b11101111001,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110110010100: edge_mask_reg_512p3[51] <= 1'b1;
 		default: edge_mask_reg_512p3[51] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000101100,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100011001,
12'b11100011010,
12'b11100011011,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b100000010111,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000101010,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100000111010,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010110,
12'b100101010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010110,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100100110,
12'b110100110101,
12'b110100110110,
12'b110101000101: edge_mask_reg_512p3[52] <= 1'b1;
 		default: edge_mask_reg_512p3[52] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101011001,
12'b11101011010,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b110001100101,
12'b110001110100,
12'b110001110101,
12'b110101110101: edge_mask_reg_512p3[53] <= 1'b1;
 		default: edge_mask_reg_512p3[53] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101110110110,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b110011000100,
12'b110011000101,
12'b110011010100,
12'b110011010101,
12'b110111000101,
12'b110111010101: edge_mask_reg_512p3[54] <= 1'b1;
 		default: edge_mask_reg_512p3[54] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111111001,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100110110101,
12'b100110110110,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111100101,
12'b100111100110,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b110011000100,
12'b110011000101,
12'b110011010100,
12'b110011010101,
12'b110011100100,
12'b110011100101: edge_mask_reg_512p3[55] <= 1'b1;
 		default: edge_mask_reg_512p3[55] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b100001100111,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001110101,
12'b111001110110,
12'b111010000101,
12'b111010000110: edge_mask_reg_512p3[56] <= 1'b1;
 		default: edge_mask_reg_512p3[56] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001001010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011001,
12'b11101011010,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b100001100111,
12'b100001101000,
12'b100001110111,
12'b100001111000,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101101100110,
12'b101101100111,
12'b101101110110,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110101100101,
12'b110101100110,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[57] <= 1'b1;
 		default: edge_mask_reg_512p3[57] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001001010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011001,
12'b11101011010,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011010,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110101100110,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001100110,
12'b111001110110: edge_mask_reg_512p3[58] <= 1'b1;
 		default: edge_mask_reg_512p3[58] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111000,
12'b100111001,
12'b101001001,
12'b101001010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001010,
12'b1101001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100111001,
12'b11100111010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100101,
12'b101100100110,
12'b110000010100,
12'b110000010101,
12'b110000010110,
12'b110000100101,
12'b110000100110,
12'b110100010101,
12'b110100100101: edge_mask_reg_512p3[59] <= 1'b1;
 		default: edge_mask_reg_512p3[59] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010010101,
12'b110010100100,
12'b110010100101: edge_mask_reg_512p3[60] <= 1'b1;
 		default: edge_mask_reg_512p3[60] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101: edge_mask_reg_512p3[61] <= 1'b1;
 		default: edge_mask_reg_512p3[61] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000110111,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000100101,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10100011000,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001101001,
12'b11001101010,
12'b11100010101,
12'b11100011001,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010100,
12'b100001010101,
12'b100100100011,
12'b100100100100,
12'b100100110011,
12'b100100110100,
12'b100101000011,
12'b100101000100,
12'b101000100011,
12'b101000100100,
12'b101000110011,
12'b101000110100,
12'b101001000011,
12'b101001000100,
12'b101100100100,
12'b101100110100: edge_mask_reg_512p3[62] <= 1'b1;
 		default: edge_mask_reg_512p3[62] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001010,
12'b11101001011,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100101010111,
12'b100101011000,
12'b100101011001,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b101001010111,
12'b101001011000,
12'b101001011001,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101101001,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110101010111,
12'b110101011000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b111001010111,
12'b111001100110,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111101100110,
12'b111101100111: edge_mask_reg_512p3[63] <= 1'b1;
 		default: edge_mask_reg_512p3[63] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101001000101,
12'b101001000110,
12'b101100010100,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000100100,
12'b110000100101,
12'b110000100110,
12'b110000110100,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[64] <= 1'b1;
 		default: edge_mask_reg_512p3[64] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011010,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001011001,
12'b10001011010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101011010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101001001,
12'b11101001010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100100100,
12'b101100100101,
12'b101100110100,
12'b101100110101,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000110100: edge_mask_reg_512p3[65] <= 1'b1;
 		default: edge_mask_reg_512p3[65] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001000011,
12'b101001000100,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[66] <= 1'b1;
 		default: edge_mask_reg_512p3[66] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001000011,
12'b101001000100,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[67] <= 1'b1;
 		default: edge_mask_reg_512p3[67] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001000100,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101000100,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[68] <= 1'b1;
 		default: edge_mask_reg_512p3[68] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001000100,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101000100,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[69] <= 1'b1;
 		default: edge_mask_reg_512p3[69] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100101001,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101000100,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[70] <= 1'b1;
 		default: edge_mask_reg_512p3[70] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110110010110,
12'b110110010111,
12'b110110100110,
12'b110110100111,
12'b110110110110,
12'b111010010111,
12'b111010100110,
12'b111010100111: edge_mask_reg_512p3[71] <= 1'b1;
 		default: edge_mask_reg_512p3[71] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110111000101,
12'b110111010101: edge_mask_reg_512p3[72] <= 1'b1;
 		default: edge_mask_reg_512p3[72] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110111000101,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[73] <= 1'b1;
 		default: edge_mask_reg_512p3[73] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111000101,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[74] <= 1'b1;
 		default: edge_mask_reg_512p3[74] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111000101,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[75] <= 1'b1;
 		default: edge_mask_reg_512p3[75] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011011010,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011101010,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111001000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111011000,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011010111,
12'b110011100101,
12'b110011100110,
12'b110011100111,
12'b110111000101,
12'b110111000110,
12'b110111010101,
12'b110111010110,
12'b110111100101,
12'b110111100110,
12'b111011010110,
12'b111011100110: edge_mask_reg_512p3[76] <= 1'b1;
 		default: edge_mask_reg_512p3[76] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001110101,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110110000100,
12'b110110000101,
12'b110110010101: edge_mask_reg_512p3[77] <= 1'b1;
 		default: edge_mask_reg_512p3[77] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b110001110101,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110110000101: edge_mask_reg_512p3[78] <= 1'b1;
 		default: edge_mask_reg_512p3[78] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111011,
12'b10001111100,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101111011,
12'b10101111100,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10110111101,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b11001111011,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010101101,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11010111101,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11110111100,
12'b11111001010,
12'b11111001011,
12'b11111001100,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100010111010,
12'b100010111011,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110110100111,
12'b110110110110,
12'b110110110111,
12'b111010110110,
12'b111010110111: edge_mask_reg_512p3[79] <= 1'b1;
 		default: edge_mask_reg_512p3[79] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b10000100101,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11100010101,
12'b11100010110,
12'b11100011001,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101000,
12'b11100101001,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100111000,
12'b11100111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b100000010100,
12'b100000010101,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100100010100,
12'b100100010101,
12'b100100100011,
12'b100100100100,
12'b100100100101,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b101000100011,
12'b101000100100,
12'b101000100101,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101001000011,
12'b101100100100,
12'b101100110100: edge_mask_reg_512p3[80] <= 1'b1;
 		default: edge_mask_reg_512p3[80] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101011,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111011,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010100101,
12'b110010100110,
12'b110010110101,
12'b110010110110,
12'b110110100110,
12'b110110110110: edge_mask_reg_512p3[81] <= 1'b1;
 		default: edge_mask_reg_512p3[81] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010101,
12'b110001110101,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110110000101: edge_mask_reg_512p3[82] <= 1'b1;
 		default: edge_mask_reg_512p3[82] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b110000000110,
12'b110000000111,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010110,
12'b111000000110,
12'b111000010110,
12'b111100000110: edge_mask_reg_512p3[83] <= 1'b1;
 		default: edge_mask_reg_512p3[83] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011010,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100101100110,
12'b100101100111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010110,
12'b100110010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b110001100101,
12'b110001100110,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110101100101,
12'b110101100110,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001110110: edge_mask_reg_512p3[84] <= 1'b1;
 		default: edge_mask_reg_512p3[84] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100010101,
12'b100100010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[85] <= 1'b1;
 		default: edge_mask_reg_512p3[85] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101001000111,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[86] <= 1'b1;
 		default: edge_mask_reg_512p3[86] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000110,
12'b100101000111,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101001000111,
12'b101100010100,
12'b101100010101,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000010101,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[87] <= 1'b1;
 		default: edge_mask_reg_512p3[87] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000110,
12'b100101000111,
12'b101000010101,
12'b101000010110,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101001000111,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110101,
12'b101100110110,
12'b110000010101,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100010101,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[88] <= 1'b1;
 		default: edge_mask_reg_512p3[88] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011010,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101001000111,
12'b101100100101,
12'b101100100110,
12'b101100110101,
12'b101100110110,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[89] <= 1'b1;
 		default: edge_mask_reg_512p3[89] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101101010,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100101,
12'b101100100110,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b110000100101,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100110101,
12'b110100110110,
12'b110101000101,
12'b110101000110: edge_mask_reg_512p3[90] <= 1'b1;
 		default: edge_mask_reg_512p3[90] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101100101,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001100101,
12'b101001100110,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b110001110101,
12'b110001110110,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010100,
12'b110010010101,
12'b110101110101,
12'b110101110110,
12'b110110000100,
12'b110110000101,
12'b110110010100,
12'b110110010101,
12'b111001110101,
12'b111010000101: edge_mask_reg_512p3[91] <= 1'b1;
 		default: edge_mask_reg_512p3[91] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101000,
12'b10011101001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101001,
12'b11010001000,
12'b11010001001,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111011001,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010100,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010100100,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110100100,
12'b110110110100,
12'b110110110101,
12'b110111000100,
12'b110111000101: edge_mask_reg_512p3[92] <= 1'b1;
 		default: edge_mask_reg_512p3[92] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011010100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101111000100,
12'b110010100100,
12'b110010110100: edge_mask_reg_512p3[93] <= 1'b1;
 		default: edge_mask_reg_512p3[93] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010101,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011010100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010110100: edge_mask_reg_512p3[94] <= 1'b1;
 		default: edge_mask_reg_512p3[94] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011010100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100: edge_mask_reg_512p3[95] <= 1'b1;
 		default: edge_mask_reg_512p3[95] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110111001,
12'b11110111010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b101010010100,
12'b101010100100: edge_mask_reg_512p3[96] <= 1'b1;
 		default: edge_mask_reg_512p3[96] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111001,
12'b10100111010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101101010100,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b110001100100: edge_mask_reg_512p3[97] <= 1'b1;
 		default: edge_mask_reg_512p3[97] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110110010101,
12'b110110010110,
12'b110110100101,
12'b111010010101: edge_mask_reg_512p3[98] <= 1'b1;
 		default: edge_mask_reg_512p3[98] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011010,
12'b11111011011,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100010111010,
12'b100010111011,
12'b100011001000,
12'b100011001001,
12'b100110010111,
12'b100110011000,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b100111000111,
12'b100111001000,
12'b100111001001,
12'b101010010111,
12'b101010011000,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101010110111,
12'b101010111000,
12'b101010111001,
12'b101011000111,
12'b101011001000,
12'b101011001001,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b101111000111,
12'b101111001000,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110011000110,
12'b110011000111,
12'b110011001000,
12'b110110010111,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b110110110111,
12'b110110111000,
12'b110111000110,
12'b110111000111,
12'b110111001000,
12'b111010100110,
12'b111010100111,
12'b111010110110,
12'b111010110111,
12'b111110100110,
12'b111110110110,
12'b111110110111: edge_mask_reg_512p3[99] <= 1'b1;
 		default: edge_mask_reg_512p3[99] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011010,
12'b11111011011,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100010111010,
12'b100010111011,
12'b100011001000,
12'b100011001001,
12'b100110010111,
12'b100110011000,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b100111000111,
12'b100111001000,
12'b100111001001,
12'b101010010111,
12'b101010011000,
12'b101010100111,
12'b101010101000,
12'b101010110111,
12'b101010111000,
12'b101010111001,
12'b101011000111,
12'b101011001000,
12'b101011001001,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b101111000111,
12'b101111001000,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110011000110,
12'b110011000111,
12'b110011001000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b110110110111,
12'b110110111000,
12'b110111000110,
12'b110111000111,
12'b110111001000,
12'b111010100110,
12'b111010100111,
12'b111010110110,
12'b111010110111: edge_mask_reg_512p3[100] <= 1'b1;
 		default: edge_mask_reg_512p3[100] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011001,
12'b11011011010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111001001,
12'b11111001010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b100111000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101011000011,
12'b101011000100,
12'b101110010100,
12'b101110100100: edge_mask_reg_512p3[101] <= 1'b1;
 		default: edge_mask_reg_512p3[101] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b10111011010,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111001001,
12'b11111001010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b100111000100,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101011000011,
12'b101011000100,
12'b101110100100: edge_mask_reg_512p3[102] <= 1'b1;
 		default: edge_mask_reg_512p3[102] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b100001100101,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101110000100: edge_mask_reg_512p3[103] <= 1'b1;
 		default: edge_mask_reg_512p3[103] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111010,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101101001,
12'b11101101010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100110100,
12'b100100110101,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b101000100100,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101100110100,
12'b101101000100,
12'b101101010100: edge_mask_reg_512p3[104] <= 1'b1;
 		default: edge_mask_reg_512p3[104] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b101000100100,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101001000101,
12'b101100110100,
12'b101101000100: edge_mask_reg_512p3[105] <= 1'b1;
 		default: edge_mask_reg_512p3[105] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p3[106] <= 1'b1;
 		default: edge_mask_reg_512p3[106] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111010,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101110000100,
12'b101110000101,
12'b101110010100: edge_mask_reg_512p3[107] <= 1'b1;
 		default: edge_mask_reg_512p3[107] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101101110100,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p3[108] <= 1'b1;
 		default: edge_mask_reg_512p3[108] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p3[109] <= 1'b1;
 		default: edge_mask_reg_512p3[109] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p3[110] <= 1'b1;
 		default: edge_mask_reg_512p3[110] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001100101,
12'b101001100110,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101101100110,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010100,
12'b110010010101,
12'b110101110101,
12'b110110000101,
12'b110110010101: edge_mask_reg_512p3[111] <= 1'b1;
 		default: edge_mask_reg_512p3[111] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110101,
12'b101110110,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000101,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101110100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110111001,
12'b11110111010,
12'b11110111011: edge_mask_reg_512p3[112] <= 1'b1;
 		default: edge_mask_reg_512p3[112] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b110110110110,
12'b111010100101: edge_mask_reg_512p3[113] <= 1'b1;
 		default: edge_mask_reg_512p3[113] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000110,
12'b100011000111,
12'b100110010101,
12'b100110010110,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b100111000110,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101111000100,
12'b101111000101,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101,
12'b110011000101,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p3[114] <= 1'b1;
 		default: edge_mask_reg_512p3[114] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101111000100,
12'b101111000101,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b110111000100,
12'b110111000101: edge_mask_reg_512p3[115] <= 1'b1;
 		default: edge_mask_reg_512p3[115] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100101,
12'b110010100110,
12'b110010110101,
12'b110010110110,
12'b110110100101,
12'b110110100110,
12'b110110110101,
12'b110110110110,
12'b111010100101,
12'b111010110101: edge_mask_reg_512p3[116] <= 1'b1;
 		default: edge_mask_reg_512p3[116] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010100,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b110010110100,
12'b110011000100: edge_mask_reg_512p3[117] <= 1'b1;
 		default: edge_mask_reg_512p3[117] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110000101,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010000100,
12'b11010000101,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101010,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b11111011010,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100100,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101: edge_mask_reg_512p3[118] <= 1'b1;
 		default: edge_mask_reg_512p3[118] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100111001,
12'b11100111010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b101100100110,
12'b101100100111,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110000100101,
12'b110000100110,
12'b110000100111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b110100010111,
12'b110100100101,
12'b110100100110,
12'b111000000101,
12'b111000000110,
12'b111000010101,
12'b111000010110,
12'b111000100101,
12'b111000100110,
12'b111100000110,
12'b111100010110: edge_mask_reg_512p3[119] <= 1'b1;
 		default: edge_mask_reg_512p3[119] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b110010110100,
12'b110011000100,
12'b110011010100: edge_mask_reg_512p3[120] <= 1'b1;
 		default: edge_mask_reg_512p3[120] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000101,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b10111011010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000011,
12'b11111001001,
12'b11111001010,
12'b100010010011,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100011000011,
12'b100110100011,
12'b100110110011: edge_mask_reg_512p3[121] <= 1'b1;
 		default: edge_mask_reg_512p3[121] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001000101,
12'b101001000110,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110101010101,
12'b110101100101,
12'b110101100110,
12'b110101100111,
12'b110101110101,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001010101,
12'b111001100101,
12'b111001100110,
12'b111001110101,
12'b111001110110,
12'b111010000110,
12'b111101110110: edge_mask_reg_512p3[122] <= 1'b1;
 		default: edge_mask_reg_512p3[122] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010000101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110000011,
12'b10110000100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111010100,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000011,
12'b11011000100,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000011,
12'b11111001000,
12'b11111001001,
12'b100010010011,
12'b100010100011,
12'b100010110011,
12'b100010110100,
12'b100011000011,
12'b100110100011,
12'b100110110011: edge_mask_reg_512p3[123] <= 1'b1;
 		default: edge_mask_reg_512p3[123] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101101100110,
12'b101101100111,
12'b101101110110,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110101100110,
12'b110101100111,
12'b110101110101,
12'b110101110110,
12'b110101110111,
12'b110110000101,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[124] <= 1'b1;
 		default: edge_mask_reg_512p3[124] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b100001110011,
12'b100010000011,
12'b100010010011,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110010011: edge_mask_reg_512p3[125] <= 1'b1;
 		default: edge_mask_reg_512p3[125] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110111000,
12'b11110111001,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101010000011,
12'b101010010011,
12'b101010100011: edge_mask_reg_512p3[126] <= 1'b1;
 		default: edge_mask_reg_512p3[126] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100101,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110100,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110100011,
12'b11110100100,
12'b11110101000,
12'b11110101001,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101010000011,
12'b101010010011,
12'b101010100011: edge_mask_reg_512p3[127] <= 1'b1;
 		default: edge_mask_reg_512p3[127] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001111000,
12'b11001111001,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101000110100,
12'b101000110101,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100100,
12'b101001100101,
12'b101100110100,
12'b101101000100,
12'b101101000101,
12'b101101010100,
12'b101101010101,
12'b101101100100,
12'b110001000100,
12'b110001010100: edge_mask_reg_512p3[128] <= 1'b1;
 		default: edge_mask_reg_512p3[128] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110101,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110111001,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101110100100: edge_mask_reg_512p3[129] <= 1'b1;
 		default: edge_mask_reg_512p3[129] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110101,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10101101001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110111001,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101110100100: edge_mask_reg_512p3[130] <= 1'b1;
 		default: edge_mask_reg_512p3[130] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011: edge_mask_reg_512p3[131] <= 1'b1;
 		default: edge_mask_reg_512p3[131] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011: edge_mask_reg_512p3[132] <= 1'b1;
 		default: edge_mask_reg_512p3[132] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001110011: edge_mask_reg_512p3[133] <= 1'b1;
 		default: edge_mask_reg_512p3[133] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001100011,
12'b101001100100,
12'b101001110011: edge_mask_reg_512p3[134] <= 1'b1;
 		default: edge_mask_reg_512p3[134] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[135] <= 1'b1;
 		default: edge_mask_reg_512p3[135] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[136] <= 1'b1;
 		default: edge_mask_reg_512p3[136] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[137] <= 1'b1;
 		default: edge_mask_reg_512p3[137] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100: edge_mask_reg_512p3[138] <= 1'b1;
 		default: edge_mask_reg_512p3[138] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011001,
12'b10010011010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011001,
12'b10110011010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001110011: edge_mask_reg_512p3[139] <= 1'b1;
 		default: edge_mask_reg_512p3[139] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[140] <= 1'b1;
 		default: edge_mask_reg_512p3[140] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b100001000011,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100: edge_mask_reg_512p3[141] <= 1'b1;
 		default: edge_mask_reg_512p3[141] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101011010,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010111,
12'b100110011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010111,
12'b101101100110,
12'b101101100111,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b110001100110,
12'b110001100111,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110110,
12'b110101110111,
12'b110110000101,
12'b110110000110,
12'b110110000111,
12'b110110010101,
12'b110110010110,
12'b110110010111,
12'b111001110110,
12'b111010000110,
12'b111010010110: edge_mask_reg_512p3[142] <= 1'b1;
 		default: edge_mask_reg_512p3[142] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010111,
12'b100000011000,
12'b100000011001,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100001000,
12'b101100010110,
12'b101100010111,
12'b101100011000,
12'b110000000110,
12'b110000000111,
12'b110000001000,
12'b110000010110,
12'b110000010111,
12'b110000011000,
12'b110100000110,
12'b110100000111,
12'b110100010110,
12'b110100010111,
12'b111000000110,
12'b111000000111,
12'b111000010110,
12'b111000010111,
12'b111100000110,
12'b111100000111,
12'b111100010110,
12'b111100010111: edge_mask_reg_512p3[143] <= 1'b1;
 		default: edge_mask_reg_512p3[143] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100010110101,
12'b100010110110,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011000101,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[144] <= 1'b1;
 		default: edge_mask_reg_512p3[144] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011000101,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[145] <= 1'b1;
 		default: edge_mask_reg_512p3[145] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[146] <= 1'b1;
 		default: edge_mask_reg_512p3[146] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000110,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[147] <= 1'b1;
 		default: edge_mask_reg_512p3[147] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[148] <= 1'b1;
 		default: edge_mask_reg_512p3[148] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111010101,
12'b110111100101: edge_mask_reg_512p3[149] <= 1'b1;
 		default: edge_mask_reg_512p3[149] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110111010101,
12'b110111100101,
12'b110111110101: edge_mask_reg_512p3[150] <= 1'b1;
 		default: edge_mask_reg_512p3[150] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110111010101,
12'b110111100101,
12'b110111110101: edge_mask_reg_512p3[151] <= 1'b1;
 		default: edge_mask_reg_512p3[151] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110111010101,
12'b110111100101,
12'b110111100110,
12'b110111110101,
12'b110111110110: edge_mask_reg_512p3[152] <= 1'b1;
 		default: edge_mask_reg_512p3[152] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b100010110111,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110110,
12'b100111110111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110110,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110011100101,
12'b110011100110,
12'b110111000101,
12'b110111000110,
12'b110111010101,
12'b110111010110,
12'b110111100101: edge_mask_reg_512p3[153] <= 1'b1;
 		default: edge_mask_reg_512p3[153] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111011,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011000,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11101011011,
12'b11101101000,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011010,
12'b11110011011,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010001011,
12'b100010010111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010111,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b110110000111,
12'b111010000110,
12'b111010000111: edge_mask_reg_512p3[154] <= 1'b1;
 		default: edge_mask_reg_512p3[154] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101001110011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[155] <= 1'b1;
 		default: edge_mask_reg_512p3[155] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101110000100,
12'b101110010100: edge_mask_reg_512p3[156] <= 1'b1;
 		default: edge_mask_reg_512p3[156] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110100011,
12'b11110101000,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101001110011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011: edge_mask_reg_512p3[157] <= 1'b1;
 		default: edge_mask_reg_512p3[157] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101001110011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100100: edge_mask_reg_512p3[158] <= 1'b1;
 		default: edge_mask_reg_512p3[158] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110110,
12'b100100110111,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110110,
12'b101000110111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110110,
12'b101100110111,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110000100101,
12'b110000100110,
12'b110000100111,
12'b110100010101,
12'b110100010110,
12'b110100100101,
12'b110100100110,
12'b111000010101,
12'b111000010110,
12'b111000100101,
12'b111000100110,
12'b111100010110: edge_mask_reg_512p3[159] <= 1'b1;
 		default: edge_mask_reg_512p3[159] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110110101: edge_mask_reg_512p3[160] <= 1'b1;
 		default: edge_mask_reg_512p3[160] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110110101: edge_mask_reg_512p3[161] <= 1'b1;
 		default: edge_mask_reg_512p3[161] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110110101: edge_mask_reg_512p3[162] <= 1'b1;
 		default: edge_mask_reg_512p3[162] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011010,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011010,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001001,
12'b11110001010,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101101010110,
12'b101101010111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110101100101,
12'b110101100110,
12'b110101110101,
12'b110101110110: edge_mask_reg_512p3[163] <= 1'b1;
 		default: edge_mask_reg_512p3[163] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010001010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100100,
12'b101010010100: edge_mask_reg_512p3[164] <= 1'b1;
 		default: edge_mask_reg_512p3[164] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101110101,
12'b11101110110,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110100100: edge_mask_reg_512p3[165] <= 1'b1;
 		default: edge_mask_reg_512p3[165] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111001,
12'b1010111010,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000110,
12'b100011000111,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010100101,
12'b110010110101: edge_mask_reg_512p3[166] <= 1'b1;
 		default: edge_mask_reg_512p3[166] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001101011,
12'b10001101100,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010000110,
12'b100010000111,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110000111,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b110010010110,
12'b110010100110,
12'b110010100111,
12'b110010110110,
12'b110110100110,
12'b110110110110: edge_mask_reg_512p3[167] <= 1'b1;
 		default: edge_mask_reg_512p3[167] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010111,
12'b100011011000,
12'b100011011001,
12'b100011011010,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111000111,
12'b100111010110,
12'b100111010111,
12'b100111011000,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110111,
12'b100111111000,
12'b101011010110,
12'b101011010111,
12'b101011011000,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101011110111,
12'b101011111000,
12'b101111010110,
12'b101111010111,
12'b101111011000,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011010110,
12'b110011010111,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111010110,
12'b110111010111,
12'b110111100110,
12'b110111100111,
12'b110111110110,
12'b110111110111,
12'b111011010110,
12'b111011010111,
12'b111011100110,
12'b111011100111,
12'b111011110110,
12'b111011110111,
12'b111111010110,
12'b111111100110,
12'b111111100111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[168] <= 1'b1;
 		default: edge_mask_reg_512p3[168] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101110010100,
12'b101110100100: edge_mask_reg_512p3[169] <= 1'b1;
 		default: edge_mask_reg_512p3[169] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000101,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001110011,
12'b11001110100,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101110011,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b100010000011,
12'b100010010011: edge_mask_reg_512p3[170] <= 1'b1;
 		default: edge_mask_reg_512p3[170] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010111000,
12'b100010111001,
12'b100110001000,
12'b100110001001,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b101010000111,
12'b101010001000,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101010110111,
12'b101010111000,
12'b101010111001,
12'b101110001000,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110111,
12'b101110111000,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b110110110111,
12'b110110111000,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111010110110,
12'b111010110111,
12'b111110100110,
12'b111110100111,
12'b111110110110,
12'b111110110111: edge_mask_reg_512p3[171] <= 1'b1;
 		default: edge_mask_reg_512p3[171] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111010,
12'b11110111011,
12'b100010001000,
12'b100010001001,
12'b100010011000,
12'b100010011001,
12'b100010011011,
12'b100010101000,
12'b100010101001,
12'b100010101011,
12'b100110000111,
12'b100110001000,
12'b100110001001,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110101000,
12'b100110101001,
12'b101010000111,
12'b101010001000,
12'b101010001001,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101110000111,
12'b101110001000,
12'b101110010111,
12'b101110011000,
12'b101110011001,
12'b101110100111,
12'b101110101000,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110000111,
12'b110110001000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111110010111,
12'b111110100111: edge_mask_reg_512p3[172] <= 1'b1;
 		default: edge_mask_reg_512p3[172] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011010,
12'b10111011011,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010111000,
12'b100110001000,
12'b100110001001,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b101010000111,
12'b101010001000,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101010110111,
12'b101010111000,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110111,
12'b101110111000,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111: edge_mask_reg_512p3[173] <= 1'b1;
 		default: edge_mask_reg_512p3[173] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011010,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001010,
12'b10010001011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001010,
12'b10110001011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001010,
12'b11010001011,
12'b11100111010,
12'b11100111011,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111010,
12'b11101111011,
12'b100001001000,
12'b100001001001,
12'b100001011000,
12'b100001011001,
12'b100001011011,
12'b100001101000,
12'b100001101001,
12'b100001101011,
12'b100101001000,
12'b100101001001,
12'b100101011000,
12'b100101011001,
12'b100101101000,
12'b100101101001,
12'b101001000111,
12'b101001001000,
12'b101001001001,
12'b101001010111,
12'b101001011000,
12'b101001011001,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101101000111,
12'b101101001000,
12'b101101001001,
12'b101101010111,
12'b101101011000,
12'b101101011001,
12'b101101100111,
12'b101101101000,
12'b101101101001,
12'b110001000111,
12'b110001001000,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110101000111,
12'b110101001000,
12'b110101010110,
12'b110101010111,
12'b110101011000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b111001010111,
12'b111001011000,
12'b111001100111,
12'b111101010111,
12'b111101100111: edge_mask_reg_512p3[174] <= 1'b1;
 		default: edge_mask_reg_512p3[174] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[175] <= 1'b1;
 		default: edge_mask_reg_512p3[175] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[176] <= 1'b1;
 		default: edge_mask_reg_512p3[176] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[177] <= 1'b1;
 		default: edge_mask_reg_512p3[177] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[178] <= 1'b1;
 		default: edge_mask_reg_512p3[178] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[179] <= 1'b1;
 		default: edge_mask_reg_512p3[179] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[180] <= 1'b1;
 		default: edge_mask_reg_512p3[180] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[181] <= 1'b1;
 		default: edge_mask_reg_512p3[181] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[182] <= 1'b1;
 		default: edge_mask_reg_512p3[182] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[183] <= 1'b1;
 		default: edge_mask_reg_512p3[183] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[184] <= 1'b1;
 		default: edge_mask_reg_512p3[184] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[185] <= 1'b1;
 		default: edge_mask_reg_512p3[185] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[186] <= 1'b1;
 		default: edge_mask_reg_512p3[186] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[187] <= 1'b1;
 		default: edge_mask_reg_512p3[187] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[188] <= 1'b1;
 		default: edge_mask_reg_512p3[188] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[189] <= 1'b1;
 		default: edge_mask_reg_512p3[189] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011: edge_mask_reg_512p3[190] <= 1'b1;
 		default: edge_mask_reg_512p3[190] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011: edge_mask_reg_512p3[191] <= 1'b1;
 		default: edge_mask_reg_512p3[191] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011: edge_mask_reg_512p3[192] <= 1'b1;
 		default: edge_mask_reg_512p3[192] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[193] <= 1'b1;
 		default: edge_mask_reg_512p3[193] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[194] <= 1'b1;
 		default: edge_mask_reg_512p3[194] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[195] <= 1'b1;
 		default: edge_mask_reg_512p3[195] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[196] <= 1'b1;
 		default: edge_mask_reg_512p3[196] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[197] <= 1'b1;
 		default: edge_mask_reg_512p3[197] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011: edge_mask_reg_512p3[198] <= 1'b1;
 		default: edge_mask_reg_512p3[198] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011: edge_mask_reg_512p3[199] <= 1'b1;
 		default: edge_mask_reg_512p3[199] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011: edge_mask_reg_512p3[200] <= 1'b1;
 		default: edge_mask_reg_512p3[200] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[201] <= 1'b1;
 		default: edge_mask_reg_512p3[201] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[202] <= 1'b1;
 		default: edge_mask_reg_512p3[202] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[203] <= 1'b1;
 		default: edge_mask_reg_512p3[203] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[204] <= 1'b1;
 		default: edge_mask_reg_512p3[204] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000011: edge_mask_reg_512p3[205] <= 1'b1;
 		default: edge_mask_reg_512p3[205] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011: edge_mask_reg_512p3[206] <= 1'b1;
 		default: edge_mask_reg_512p3[206] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[207] <= 1'b1;
 		default: edge_mask_reg_512p3[207] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[208] <= 1'b1;
 		default: edge_mask_reg_512p3[208] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100101,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[209] <= 1'b1;
 		default: edge_mask_reg_512p3[209] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101100101,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001100100,
12'b10001100101,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100101110011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[210] <= 1'b1;
 		default: edge_mask_reg_512p3[210] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[211] <= 1'b1;
 		default: edge_mask_reg_512p3[211] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100: edge_mask_reg_512p3[212] <= 1'b1;
 		default: edge_mask_reg_512p3[212] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110111001,
12'b11110111010,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100: edge_mask_reg_512p3[213] <= 1'b1;
 		default: edge_mask_reg_512p3[213] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110111001,
12'b11110111010,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100: edge_mask_reg_512p3[214] <= 1'b1;
 		default: edge_mask_reg_512p3[214] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110101,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100: edge_mask_reg_512p3[215] <= 1'b1;
 		default: edge_mask_reg_512p3[215] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010111000,
12'b11010111001,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110100011,
12'b11110100100,
12'b11110101000,
12'b11110101001,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101101110100,
12'b101110000100,
12'b101110010100: edge_mask_reg_512p3[216] <= 1'b1;
 		default: edge_mask_reg_512p3[216] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10011011010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010000100,
12'b100010000101,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b110010010100,
12'b110010100100: edge_mask_reg_512p3[217] <= 1'b1;
 		default: edge_mask_reg_512p3[217] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10011011010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010000100,
12'b100010000101,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b110010010100,
12'b110010100100: edge_mask_reg_512p3[218] <= 1'b1;
 		default: edge_mask_reg_512p3[218] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110101,
12'b101010110110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110110010100,
12'b110110010101,
12'b110110100100,
12'b110110100101: edge_mask_reg_512p3[219] <= 1'b1;
 		default: edge_mask_reg_512p3[219] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101010,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b101001100110,
12'b101001100111,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101101100110,
12'b101101100111,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b110110000111,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111010000111,
12'b111101110110,
12'b111110000110: edge_mask_reg_512p3[220] <= 1'b1;
 		default: edge_mask_reg_512p3[220] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111010,
12'b11110111011,
12'b11111000110,
12'b11111000111,
12'b11111001010,
12'b11111001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101011,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111011,
12'b100011000101,
12'b100011000110,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b100111000110,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000101,
12'b101011000110,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000101,
12'b101111000110,
12'b110010100101,
12'b110010100110,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110110100110,
12'b110110110101,
12'b110110110110,
12'b110111000110: edge_mask_reg_512p3[221] <= 1'b1;
 		default: edge_mask_reg_512p3[221] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000111,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b101001010110,
12'b101001010111,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101101010110,
12'b101101010111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110101100101,
12'b110101100110,
12'b110101100111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[222] <= 1'b1;
 		default: edge_mask_reg_512p3[222] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000110111,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100101,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10100011000,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010100,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100100100011,
12'b100100100100,
12'b100100100101,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b101000100100,
12'b101000110100,
12'b101000110101,
12'b101001000100: edge_mask_reg_512p3[223] <= 1'b1;
 		default: edge_mask_reg_512p3[223] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111010,
12'b11110111011,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110110,
12'b110110010101,
12'b110110010110,
12'b110110100101,
12'b110110100110: edge_mask_reg_512p3[224] <= 1'b1;
 		default: edge_mask_reg_512p3[224] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111010,
12'b10110111011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111010,
12'b11010111011,
12'b11101101010,
12'b11101101011,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110101010,
12'b11110101011,
12'b100001111000,
12'b100001111001,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010001011,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100101111000,
12'b100101111001,
12'b100110000111,
12'b100110001000,
12'b100110001001,
12'b100110011000,
12'b100110011001,
12'b101001110111,
12'b101001111000,
12'b101010000111,
12'b101010001000,
12'b101010001001,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110011001,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b111010000110,
12'b111010000111,
12'b111010010110,
12'b111010010111,
12'b111110010111: edge_mask_reg_512p3[225] <= 1'b1;
 		default: edge_mask_reg_512p3[225] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110101,
12'b101110110,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101010011,
12'b10101010100,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101101000,
12'b11101101001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110101001,
12'b100001110011,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101010000011,
12'b101010010011: edge_mask_reg_512p3[226] <= 1'b1;
 		default: edge_mask_reg_512p3[226] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110101,
12'b101110110,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101010011,
12'b10101010100,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11101101000,
12'b11101101001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110101000,
12'b11110101001,
12'b100001110011,
12'b100010000011,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100110000011,
12'b100110010011,
12'b101010010011: edge_mask_reg_512p3[227] <= 1'b1;
 		default: edge_mask_reg_512p3[227] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111000,
12'b100111001,
12'b101001010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100100101,
12'b100100100110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100101,
12'b101000100110,
12'b101100010100,
12'b101100010101,
12'b110000010100,
12'b110000010101: edge_mask_reg_512p3[228] <= 1'b1;
 		default: edge_mask_reg_512p3[228] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010101,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101010100,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100010,
12'b11101101000,
12'b11101101001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101010000011: edge_mask_reg_512p3[229] <= 1'b1;
 		default: edge_mask_reg_512p3[229] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110101,
12'b1110110,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000101,
12'b10000110,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101001010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101010011,
12'b10101010100,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100010,
12'b11101100011,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110011001,
12'b100001110011,
12'b100010000011,
12'b100010010011: edge_mask_reg_512p3[230] <= 1'b1;
 		default: edge_mask_reg_512p3[230] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110111001,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101110010100,
12'b101110100100,
12'b101110110100: edge_mask_reg_512p3[231] <= 1'b1;
 		default: edge_mask_reg_512p3[231] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001101001,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110111001,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101110000100,
12'b101110010100,
12'b101110100100,
12'b101110110100,
12'b110010010100: edge_mask_reg_512p3[232] <= 1'b1;
 		default: edge_mask_reg_512p3[232] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010000110,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110010101,
12'b110110100100,
12'b110110100101,
12'b110110110101,
12'b110110110110,
12'b111010100101: edge_mask_reg_512p3[233] <= 1'b1;
 		default: edge_mask_reg_512p3[233] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000110,
12'b11110001001,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b100010000101,
12'b100010000110,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110100,
12'b110010110101,
12'b110110010101,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b111010100101: edge_mask_reg_512p3[234] <= 1'b1;
 		default: edge_mask_reg_512p3[234] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000110,
12'b11110001001,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b100010000101,
12'b100010000110,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110010101,
12'b110110100100,
12'b110110100101,
12'b110110100110,
12'b110110110101,
12'b110110110110,
12'b111010100101,
12'b111010110101: edge_mask_reg_512p3[235] <= 1'b1;
 		default: edge_mask_reg_512p3[235] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101100101,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001100110,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b110001110101,
12'b110001110110,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010100,
12'b110010010101,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101: edge_mask_reg_512p3[236] <= 1'b1;
 		default: edge_mask_reg_512p3[236] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001010101,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100101100100,
12'b100101100101,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101101100100,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b110001110100: edge_mask_reg_512p3[237] <= 1'b1;
 		default: edge_mask_reg_512p3[237] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10001001001,
12'b10001001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010101,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001010101,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101101100100,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b110001110100: edge_mask_reg_512p3[238] <= 1'b1;
 		default: edge_mask_reg_512p3[238] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b100111000110,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101111000101,
12'b101111000110,
12'b110010100101,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110110110101,
12'b110111000101: edge_mask_reg_512p3[239] <= 1'b1;
 		default: edge_mask_reg_512p3[239] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011010,
12'b11010011011,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101101010110,
12'b101101010111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110101100101,
12'b110101100110,
12'b110101110110,
12'b110101110111,
12'b111001110110: edge_mask_reg_512p3[240] <= 1'b1;
 		default: edge_mask_reg_512p3[240] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101010,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011010,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010001000,
12'b100010001001,
12'b100101010111,
12'b100101011000,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b100110001000,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101010000111,
12'b101010001000,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110101010111,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b111001100110,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111010000111,
12'b111101100110,
12'b111101100111,
12'b111101110110,
12'b111101110111,
12'b111110000110,
12'b111110000111: edge_mask_reg_512p3[241] <= 1'b1;
 		default: edge_mask_reg_512p3[241] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001101000,
12'b1001101001,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1100111001,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001000101,
12'b11001001000,
12'b11001001001,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101000101,
12'b11101001000,
12'b11101001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101101010100,
12'b101101100100: edge_mask_reg_512p3[242] <= 1'b1;
 		default: edge_mask_reg_512p3[242] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101100000110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110000100101,
12'b110000100110,
12'b110100000101,
12'b110100010101,
12'b110100100101: edge_mask_reg_512p3[243] <= 1'b1;
 		default: edge_mask_reg_512p3[243] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100010101: edge_mask_reg_512p3[244] <= 1'b1;
 		default: edge_mask_reg_512p3[244] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11100111001,
12'b11100111010,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111001,
12'b11101111010,
12'b100001000111,
12'b100001001000,
12'b100001001001,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100101000111,
12'b100101001000,
12'b100101001001,
12'b100101010111,
12'b100101011000,
12'b100101011001,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b101001000111,
12'b101001001000,
12'b101001001001,
12'b101001010111,
12'b101001011000,
12'b101001011001,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101101000111,
12'b101101001000,
12'b101101010111,
12'b101101011000,
12'b101101011001,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001000111,
12'b110001001000,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110101000111,
12'b110101001000,
12'b110101010110,
12'b110101010111,
12'b110101011000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b111001000111,
12'b111001001000,
12'b111001010110,
12'b111001010111,
12'b111001011000,
12'b111001100110,
12'b111001100111,
12'b111001101000,
12'b111101010110,
12'b111101010111,
12'b111101100110,
12'b111101100111: edge_mask_reg_512p3[245] <= 1'b1;
 		default: edge_mask_reg_512p3[245] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010101,
12'b100111010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010110100: edge_mask_reg_512p3[246] <= 1'b1;
 		default: edge_mask_reg_512p3[246] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111010111,
12'b100111011000,
12'b100111100111,
12'b100111101000,
12'b100111101001,
12'b100111110111,
12'b100111111000,
12'b100111111001,
12'b101011100111,
12'b101011101000,
12'b101011101001,
12'b101011110111,
12'b101011111000,
12'b101011111001,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111100110,
12'b110111100111,
12'b110111101000,
12'b110111110110,
12'b110111110111,
12'b110111111000,
12'b111011100110,
12'b111011100111,
12'b111011110110,
12'b111011110111,
12'b111011111000,
12'b111111100110,
12'b111111100111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[247] <= 1'b1;
 		default: edge_mask_reg_512p3[247] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100101010,
12'b10100110101,
12'b10100110110,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b11000110101,
12'b11000110110,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b100000110101,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100101000011,
12'b100101000100,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b101001000100,
12'b101001010100,
12'b101001100100: edge_mask_reg_512p3[248] <= 1'b1;
 		default: edge_mask_reg_512p3[248] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100101010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b11000101001,
12'b11000101010,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11100110100,
12'b11100110101,
12'b11100111001,
12'b11100111010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100101000011,
12'b100101000100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100: edge_mask_reg_512p3[249] <= 1'b1;
 		default: edge_mask_reg_512p3[249] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010101010,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100: edge_mask_reg_512p3[250] <= 1'b1;
 		default: edge_mask_reg_512p3[250] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[251] <= 1'b1;
 		default: edge_mask_reg_512p3[251] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110111,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100010110110,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[252] <= 1'b1;
 		default: edge_mask_reg_512p3[252] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[253] <= 1'b1;
 		default: edge_mask_reg_512p3[253] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111000,
12'b10111001,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110101,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111010110,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111100101,
12'b110111100110,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[254] <= 1'b1;
 		default: edge_mask_reg_512p3[254] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111001,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010110,
12'b100011010111,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010110,
12'b100111010111,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111010110,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111100101,
12'b110111100110,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[255] <= 1'b1;
 		default: edge_mask_reg_512p3[255] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111001,
12'b11101111010,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001111000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101111000,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110101010110,
12'b110101010111,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b111001100110,
12'b111001100111,
12'b111101100110: edge_mask_reg_512p3[256] <= 1'b1;
 		default: edge_mask_reg_512p3[256] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111001,
12'b11101111010,
12'b100001001000,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001111000,
12'b100101001000,
12'b100101010111,
12'b100101011000,
12'b100101011001,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101111000,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100111,
12'b101001101000,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110101010110,
12'b110101010111,
12'b110101011000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b111001010110,
12'b111001100110,
12'b111001100111,
12'b111101100110: edge_mask_reg_512p3[257] <= 1'b1;
 		default: edge_mask_reg_512p3[257] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b100001001000,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001111000,
12'b100101001000,
12'b100101010111,
12'b100101011000,
12'b100101011001,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101111000,
12'b101001000111,
12'b101001001000,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001000111,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110101010110,
12'b110101010111,
12'b110101011000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b111001010110,
12'b111001010111,
12'b111001100110,
12'b111001100111,
12'b111101100110: edge_mask_reg_512p3[258] <= 1'b1;
 		default: edge_mask_reg_512p3[258] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100011000111,
12'b100011001000,
12'b100110000111,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010110,
12'b110010010111,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110011000110,
12'b110110010110,
12'b110110010111,
12'b110110100101,
12'b110110100110,
12'b110110100111,
12'b110110110101,
12'b110110110110,
12'b110111000110,
12'b111010100110,
12'b111010110110: edge_mask_reg_512p3[259] <= 1'b1;
 		default: edge_mask_reg_512p3[259] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110010100101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110: edge_mask_reg_512p3[260] <= 1'b1;
 		default: edge_mask_reg_512p3[260] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[261] <= 1'b1;
 		default: edge_mask_reg_512p3[261] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[262] <= 1'b1;
 		default: edge_mask_reg_512p3[262] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[263] <= 1'b1;
 		default: edge_mask_reg_512p3[263] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[264] <= 1'b1;
 		default: edge_mask_reg_512p3[264] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[265] <= 1'b1;
 		default: edge_mask_reg_512p3[265] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[266] <= 1'b1;
 		default: edge_mask_reg_512p3[266] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[267] <= 1'b1;
 		default: edge_mask_reg_512p3[267] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[268] <= 1'b1;
 		default: edge_mask_reg_512p3[268] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[269] <= 1'b1;
 		default: edge_mask_reg_512p3[269] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[270] <= 1'b1;
 		default: edge_mask_reg_512p3[270] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[271] <= 1'b1;
 		default: edge_mask_reg_512p3[271] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[272] <= 1'b1;
 		default: edge_mask_reg_512p3[272] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[273] <= 1'b1;
 		default: edge_mask_reg_512p3[273] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[274] <= 1'b1;
 		default: edge_mask_reg_512p3[274] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[275] <= 1'b1;
 		default: edge_mask_reg_512p3[275] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011: edge_mask_reg_512p3[276] <= 1'b1;
 		default: edge_mask_reg_512p3[276] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p3[277] <= 1'b1;
 		default: edge_mask_reg_512p3[277] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[278] <= 1'b1;
 		default: edge_mask_reg_512p3[278] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010011,
12'b100001010100,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101010011,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[279] <= 1'b1;
 		default: edge_mask_reg_512p3[279] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101000100,
12'b10101000101,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001000100,
12'b11001000101,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101000100,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011,
12'b100101110100,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[280] <= 1'b1;
 		default: edge_mask_reg_512p3[280] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110010110,
12'b110110010111,
12'b110110100110,
12'b110110100111,
12'b111010010110,
12'b111010100110,
12'b111010100111,
12'b111110100110: edge_mask_reg_512p3[281] <= 1'b1;
 		default: edge_mask_reg_512p3[281] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101101010110,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110101100101,
12'b110101100110,
12'b110101110101,
12'b110101110110: edge_mask_reg_512p3[282] <= 1'b1;
 		default: edge_mask_reg_512p3[282] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101101010110,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b110001100101,
12'b110001100110,
12'b110001110101,
12'b110001110110,
12'b110101100101,
12'b110101100110,
12'b110101110101,
12'b110101110110: edge_mask_reg_512p3[283] <= 1'b1;
 		default: edge_mask_reg_512p3[283] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011010,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011001,
12'b11110011010,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110001001,
12'b101001100110,
12'b101001100111,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010001001,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111010000111,
12'b111101110110,
12'b111101110111,
12'b111110000110,
12'b111110000111: edge_mask_reg_512p3[284] <= 1'b1;
 		default: edge_mask_reg_512p3[284] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001001,
12'b1111001010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110111001,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110010000100,
12'b110010010100,
12'b110010100100: edge_mask_reg_512p3[285] <= 1'b1;
 		default: edge_mask_reg_512p3[285] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001001,
12'b11111001010,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010110111,
12'b100010111000,
12'b100110000111,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010110,
12'b110010010111,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110110010110,
12'b110110010111,
12'b110110100101,
12'b110110100110,
12'b110110100111,
12'b110110110101,
12'b110110110110,
12'b111010100110,
12'b111010110110: edge_mask_reg_512p3[286] <= 1'b1;
 		default: edge_mask_reg_512p3[286] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101101010,
12'b11101101011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101010,
12'b11110101011,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110100100: edge_mask_reg_512p3[287] <= 1'b1;
 		default: edge_mask_reg_512p3[287] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11111001000,
12'b11111001001,
12'b100010010100,
12'b100010010101,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110010100,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000101,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101111000100,
12'b101111000101,
12'b110010100100,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110110110100,
12'b110110110101,
12'b110111000100,
12'b110111000101: edge_mask_reg_512p3[288] <= 1'b1;
 		default: edge_mask_reg_512p3[288] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000101100,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100011010,
12'b11100011011,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101101010,
12'b100000010111,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000101010,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100000111010,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010110,
12'b100101010111,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110000110111,
12'b110001000101,
12'b110001000110,
12'b110100100110,
12'b110100110101,
12'b110100110110,
12'b110101000101,
12'b110101000110: edge_mask_reg_512p3[289] <= 1'b1;
 		default: edge_mask_reg_512p3[289] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000101100,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100011001,
12'b11100011010,
12'b11100011011,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101011010,
12'b100000010111,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000101010,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100000111010,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101001000111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000110,
12'b101101000111,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110000110111,
12'b110100100101,
12'b110100100110,
12'b110100110101,
12'b110100110110: edge_mask_reg_512p3[290] <= 1'b1;
 		default: edge_mask_reg_512p3[290] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101: edge_mask_reg_512p3[291] <= 1'b1;
 		default: edge_mask_reg_512p3[291] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b110011000100,
12'b110011000101,
12'b110011010100,
12'b110011010101: edge_mask_reg_512p3[292] <= 1'b1;
 		default: edge_mask_reg_512p3[292] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b100111100101,
12'b100111100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100101,
12'b101011100110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b110011000101,
12'b110011010101: edge_mask_reg_512p3[293] <= 1'b1;
 		default: edge_mask_reg_512p3[293] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b100111100101,
12'b100111100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100101,
12'b101011100110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b110011000101,
12'b110011010101: edge_mask_reg_512p3[294] <= 1'b1;
 		default: edge_mask_reg_512p3[294] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111100100,
12'b101111100101,
12'b110011000101,
12'b110011010101,
12'b110011100101: edge_mask_reg_512p3[295] <= 1'b1;
 		default: edge_mask_reg_512p3[295] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001000100,
12'b11001000101,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001001,
12'b11110001010,
12'b100001010011,
12'b100001100011,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100010000011: edge_mask_reg_512p3[296] <= 1'b1;
 		default: edge_mask_reg_512p3[296] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000101,
12'b100111000110,
12'b101010010100,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101110010100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010100100,
12'b110010110100: edge_mask_reg_512p3[297] <= 1'b1;
 		default: edge_mask_reg_512p3[297] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000101010,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001001001,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001111000,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110111,
12'b100101111000,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110111,
12'b101101000110,
12'b101101000111,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b110001000111,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110110,
12'b110101010110,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b111001010110,
12'b111001100110,
12'b111001110110: edge_mask_reg_512p3[298] <= 1'b1;
 		default: edge_mask_reg_512p3[298] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011010,
12'b11011011011,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100010111011,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110110,
12'b110110100110,
12'b110110110110: edge_mask_reg_512p3[299] <= 1'b1;
 		default: edge_mask_reg_512p3[299] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010101,
12'b101011010110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b110010100100,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110011010101,
12'b110110110101,
12'b110111000101,
12'b110111010101: edge_mask_reg_512p3[300] <= 1'b1;
 		default: edge_mask_reg_512p3[300] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010101,
12'b101011010110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101,
12'b110011010100,
12'b110011010101,
12'b110111000101,
12'b110111010101: edge_mask_reg_512p3[301] <= 1'b1;
 		default: edge_mask_reg_512p3[301] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110110000100,
12'b110110010100,
12'b110110010101,
12'b110110100100: edge_mask_reg_512p3[302] <= 1'b1;
 		default: edge_mask_reg_512p3[302] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001001,
12'b10011001010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110010100100: edge_mask_reg_512p3[303] <= 1'b1;
 		default: edge_mask_reg_512p3[303] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001001,
12'b10011001010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101110010100,
12'b101110100100,
12'b101110100101,
12'b110010100100: edge_mask_reg_512p3[304] <= 1'b1;
 		default: edge_mask_reg_512p3[304] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101: edge_mask_reg_512p3[305] <= 1'b1;
 		default: edge_mask_reg_512p3[305] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101: edge_mask_reg_512p3[306] <= 1'b1;
 		default: edge_mask_reg_512p3[306] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010101,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10101100100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110111000,
12'b11110111001,
12'b100001110011,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010110011,
12'b100110000011,
12'b100110010011,
12'b100110100011,
12'b101010010011: edge_mask_reg_512p3[307] <= 1'b1;
 		default: edge_mask_reg_512p3[307] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010101,
12'b110010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101100100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001110011,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100: edge_mask_reg_512p3[308] <= 1'b1;
 		default: edge_mask_reg_512p3[308] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110110,
12'b11110111010,
12'b11110111011,
12'b11111001011,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100010001011,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011011,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101011,
12'b100101110110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000101,
12'b101010000110,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110110,
12'b101110000101,
12'b101110000110,
12'b101110010101,
12'b101110010110,
12'b101110100101,
12'b101110100110,
12'b101110110110,
12'b110010010110,
12'b110010100110: edge_mask_reg_512p3[309] <= 1'b1;
 		default: edge_mask_reg_512p3[309] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100100,
12'b101110000100,
12'b101110010100: edge_mask_reg_512p3[310] <= 1'b1;
 		default: edge_mask_reg_512p3[310] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100100: edge_mask_reg_512p3[311] <= 1'b1;
 		default: edge_mask_reg_512p3[311] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b101001110011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101010100100: edge_mask_reg_512p3[312] <= 1'b1;
 		default: edge_mask_reg_512p3[312] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001101010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100110000111,
12'b100110001000,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b111010000110,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111110010110: edge_mask_reg_512p3[313] <= 1'b1;
 		default: edge_mask_reg_512p3[313] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11100111001,
12'b11100111010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101001010,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101110011: edge_mask_reg_512p3[314] <= 1'b1;
 		default: edge_mask_reg_512p3[314] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000111,
12'b100110001000,
12'b101001010110,
12'b101001010111,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000111,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[315] <= 1'b1;
 		default: edge_mask_reg_512p3[315] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000111,
12'b100110001000,
12'b101001010110,
12'b101001010111,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000111,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[316] <= 1'b1;
 		default: edge_mask_reg_512p3[316] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000111,
12'b100110001000,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000111,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110101010110,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111010000110: edge_mask_reg_512p3[317] <= 1'b1;
 		default: edge_mask_reg_512p3[317] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111001,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001010,
12'b11111001011,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010111,
12'b100011011000,
12'b100011011001,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100011111010,
12'b100111010111,
12'b100111011000,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111101001,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b100111111001,
12'b101011010111,
12'b101011011000,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111010111,
12'b101111011000,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011010111,
12'b110011011000,
12'b110011100101,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111100101,
12'b110111100110,
12'b110111100111,
12'b110111110101,
12'b110111110110,
12'b110111110111,
12'b111011100110,
12'b111011100111,
12'b111011110110,
12'b111011110111,
12'b111111100110,
12'b111111110110: edge_mask_reg_512p3[318] <= 1'b1;
 		default: edge_mask_reg_512p3[318] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111001,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001010,
12'b11111001011,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111111000,
12'b11111111001,
12'b100011010111,
12'b100011011000,
12'b100011011001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111010111,
12'b100111011000,
12'b100111100111,
12'b100111101000,
12'b100111101001,
12'b100111110111,
12'b100111111000,
12'b100111111001,
12'b101011010111,
12'b101011011000,
12'b101011100111,
12'b101011101000,
12'b101011101001,
12'b101011110111,
12'b101011111000,
12'b101011111001,
12'b101111010111,
12'b101111011000,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110111,
12'b101111111000,
12'b110011010111,
12'b110011011000,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111100110,
12'b110111100111,
12'b110111101000,
12'b110111110110,
12'b110111110111,
12'b110111111000,
12'b111011100110,
12'b111011100111,
12'b111011110110,
12'b111011110111,
12'b111011111000,
12'b111111100110,
12'b111111100111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[319] <= 1'b1;
 		default: edge_mask_reg_512p3[319] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111010,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111011,
12'b1001111100,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b11000011010,
12'b11000101010,
12'b11000101011,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101010,
12'b11001101011,
12'b11100101010,
12'b11100101011,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101011010,
12'b11101011011,
12'b100000110111,
12'b100000111000,
12'b100000111001,
12'b100000111010,
12'b100000111011,
12'b100001000111,
12'b100001001000,
12'b100001001001,
12'b100001001010,
12'b100001001011,
12'b100001011000,
12'b100100101000,
12'b100100110111,
12'b100100111000,
12'b100100111001,
12'b100101000111,
12'b100101001000,
12'b100101001001,
12'b100101010111,
12'b100101011000,
12'b101000110110,
12'b101000110111,
12'b101000111000,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001010111,
12'b101001011000,
12'b101100110110,
12'b101100110111,
12'b101100111000,
12'b101101000110,
12'b101101000111,
12'b101101001000,
12'b101101011000,
12'b110000110110,
12'b110000110111,
12'b110000111000,
12'b110001000110,
12'b110001000111,
12'b110001001000,
12'b110100110110,
12'b110100110111,
12'b110101000110,
12'b110101000111,
12'b111000110110,
12'b111000110111,
12'b111001000110,
12'b111001000111,
12'b111100110111,
12'b111101000111: edge_mask_reg_512p3[320] <= 1'b1;
 		default: edge_mask_reg_512p3[320] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101101001,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b101000100101,
12'b101000100110,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101100110100,
12'b101100110101,
12'b101101000100,
12'b101101000101,
12'b101101010100,
12'b110000110100,
12'b110000110101,
12'b110001000100,
12'b110001000101: edge_mask_reg_512p3[321] <= 1'b1;
 		default: edge_mask_reg_512p3[321] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111010,
12'b11110111011,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110011001,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110101001,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110111,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111010101000,
12'b111010110111,
12'b111110010110,
12'b111110010111,
12'b111110100110,
12'b111110100111,
12'b111110110111: edge_mask_reg_512p3[322] <= 1'b1;
 		default: edge_mask_reg_512p3[322] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010101,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010100,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100101,
12'b11011101001,
12'b11011101010,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111101001,
12'b11111101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010011,
12'b100011010100,
12'b100011010101,
12'b100011010110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010011,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101,
12'b101011010100,
12'b101011010101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b110010110100,
12'b110011000100: edge_mask_reg_512p3[323] <= 1'b1;
 		default: edge_mask_reg_512p3[323] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001010,
12'b100111000,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b11000100101,
12'b11000100110,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100100101,
12'b11100100110,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b100000100101,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101100110100,
12'b101100110101,
12'b101101000100,
12'b101101000101,
12'b101101010100,
12'b110001000100: edge_mask_reg_512p3[324] <= 1'b1;
 		default: edge_mask_reg_512p3[324] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100101,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011000,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100010101,
12'b11100011001,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100100011,
12'b100100100100,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b101000100011,
12'b101000100100,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101100100100,
12'b101100110100,
12'b101100110101,
12'b101101000100,
12'b101101000101,
12'b110001000100: edge_mask_reg_512p3[325] <= 1'b1;
 		default: edge_mask_reg_512p3[325] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100011000,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000100101,
12'b11000100110,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100101000,
12'b11100101001,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011000,
12'b11101011001,
12'b11101101001,
12'b100000100100,
12'b100000100101,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010100,
12'b100101010101,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101100110100,
12'b101101000100,
12'b101101010100,
12'b110001000100: edge_mask_reg_512p3[326] <= 1'b1;
 		default: edge_mask_reg_512p3[326] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101000,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010101,
12'b10111010110,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010100,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010100,
12'b100011010101,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010011,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010110100: edge_mask_reg_512p3[327] <= 1'b1;
 		default: edge_mask_reg_512p3[327] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111001,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111001010,
12'b11111001011,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010111,
12'b100011011000,
12'b100011011001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111010111,
12'b100111011000,
12'b100111100111,
12'b100111101000,
12'b100111101001,
12'b100111110111,
12'b100111111000,
12'b100111111001,
12'b101011010111,
12'b101011011000,
12'b101011100111,
12'b101011101000,
12'b101011110111,
12'b101011111000,
12'b101111010111,
12'b101111011000,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011010111,
12'b110011011000,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111100110,
12'b110111100111,
12'b110111110110,
12'b110111110111,
12'b111011100110,
12'b111011100111,
12'b111011110110,
12'b111011110111,
12'b111111100110,
12'b111111100111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[328] <= 1'b1;
 		default: edge_mask_reg_512p3[328] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001001,
12'b11110001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001010110,
12'b101001010111,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111101110110: edge_mask_reg_512p3[329] <= 1'b1;
 		default: edge_mask_reg_512p3[329] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001001,
12'b11110001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001010110,
12'b101001010111,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b111001100110,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111101110110: edge_mask_reg_512p3[330] <= 1'b1;
 		default: edge_mask_reg_512p3[330] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111010,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b111010010110,
12'b111010010111,
12'b111010011000,
12'b111010100110,
12'b111010100111,
12'b111010101000,
12'b111110010110,
12'b111110010111,
12'b111110100110,
12'b111110100111: edge_mask_reg_512p3[331] <= 1'b1;
 		default: edge_mask_reg_512p3[331] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101011001,
12'b11101011010,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101100110101,
12'b101100110110,
12'b101101000101,
12'b101101000110,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100110101,
12'b110101000101: edge_mask_reg_512p3[332] <= 1'b1;
 		default: edge_mask_reg_512p3[332] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111011,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100100100110,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100110101,
12'b101100110110,
12'b101101000101,
12'b101101000110,
12'b110000110101,
12'b110001000101,
12'b110100110101,
12'b110101000101: edge_mask_reg_512p3[333] <= 1'b1;
 		default: edge_mask_reg_512p3[333] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001010,
12'b1011011001,
12'b1111011001,
12'b1111011010,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111100111,
12'b100111101000,
12'b100111110111,
12'b100111111000,
12'b101011100111,
12'b101011101000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111110110,
12'b110111110111,
12'b111011110110,
12'b111011110111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[334] <= 1'b1;
 		default: edge_mask_reg_512p3[334] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b110001110100,
12'b110001110101,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110101110100,
12'b110110000100,
12'b110110000101: edge_mask_reg_512p3[335] <= 1'b1;
 		default: edge_mask_reg_512p3[335] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101001,
12'b10101010,
12'b10111001,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110111010,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011000111,
12'b100011001000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100011011010,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011101010,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111000110,
12'b100111000111,
12'b100111001000,
12'b100111010110,
12'b100111010111,
12'b100111011000,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110101,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011000110,
12'b101011000111,
12'b101011010110,
12'b101011010111,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011010101,
12'b110011010110,
12'b110011010111,
12'b110011100101,
12'b110011100110,
12'b110011100111,
12'b110011110101,
12'b110011110110,
12'b110111010101,
12'b110111010110,
12'b110111100101,
12'b110111100110,
12'b110111110101,
12'b110111110110,
12'b111011010110,
12'b111011100110: edge_mask_reg_512p3[336] <= 1'b1;
 		default: edge_mask_reg_512p3[336] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110111010,
12'b111001001,
12'b111001010,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011001,
12'b11111011010,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010111,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110101,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011100101,
12'b110011100110,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111100101,
12'b110111100110,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[337] <= 1'b1;
 		default: edge_mask_reg_512p3[337] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101001001,
12'b11101001010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101: edge_mask_reg_512p3[338] <= 1'b1;
 		default: edge_mask_reg_512p3[338] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101: edge_mask_reg_512p3[339] <= 1'b1;
 		default: edge_mask_reg_512p3[339] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111000,
12'b100111001,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100101,
12'b101000100110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b110000000101,
12'b110000010100,
12'b110000010101: edge_mask_reg_512p3[340] <= 1'b1;
 		default: edge_mask_reg_512p3[340] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010101,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010110100: edge_mask_reg_512p3[341] <= 1'b1;
 		default: edge_mask_reg_512p3[341] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010110100: edge_mask_reg_512p3[342] <= 1'b1;
 		default: edge_mask_reg_512p3[342] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101000,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010101,
12'b10111010110,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010100,
12'b100011010101,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101110110100,
12'b101111000100: edge_mask_reg_512p3[343] <= 1'b1;
 		default: edge_mask_reg_512p3[343] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101001,
12'b10111101010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010110100: edge_mask_reg_512p3[344] <= 1'b1;
 		default: edge_mask_reg_512p3[344] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011010110,
12'b100011010111,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111100101,
12'b100111100110,
12'b100111100111,
12'b100111110101,
12'b100111110110,
12'b100111110111,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101011100111,
12'b101011110101,
12'b101011110110,
12'b101011110111,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110100,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011100100,
12'b110011100101,
12'b110011100110,
12'b110011110100,
12'b110011110101,
12'b110011110110,
12'b110111100101,
12'b110111110101,
12'b110111110110: edge_mask_reg_512p3[345] <= 1'b1;
 		default: edge_mask_reg_512p3[345] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111011001,
12'b11111011010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b101111000101,
12'b110010100100,
12'b110010110100,
12'b110010110101,
12'b110011000100,
12'b110011000101: edge_mask_reg_512p3[346] <= 1'b1;
 		default: edge_mask_reg_512p3[346] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011001,
12'b11011011010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000101,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110010110100: edge_mask_reg_512p3[347] <= 1'b1;
 		default: edge_mask_reg_512p3[347] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101000,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010101,
12'b10111010110,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010100,
12'b100011010101,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101110100100,
12'b101110110100,
12'b101111000100,
12'b110010110100: edge_mask_reg_512p3[348] <= 1'b1;
 		default: edge_mask_reg_512p3[348] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101110100100,
12'b101110110100,
12'b110010110100: edge_mask_reg_512p3[349] <= 1'b1;
 		default: edge_mask_reg_512p3[349] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110,
12'b111010000101,
12'b111010000110,
12'b111010010101,
12'b111010010110: edge_mask_reg_512p3[350] <= 1'b1;
 		default: edge_mask_reg_512p3[350] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001001,
12'b11010001010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100101000101,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101101010100,
12'b101101100100,
12'b101101110100,
12'b110001100100: edge_mask_reg_512p3[351] <= 1'b1;
 		default: edge_mask_reg_512p3[351] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001001,
12'b1110001010,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10100101000,
12'b10100101001,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11000110101,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11100111000,
12'b11100111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101001000,
12'b11101001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101111001,
12'b100000110100,
12'b100000110101,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100100,
12'b100001100101,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b101001000011,
12'b101001000100,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110100,
12'b101101010100,
12'b101101100100,
12'b101101110100,
12'b110001010100,
12'b110001100100: edge_mask_reg_512p3[352] <= 1'b1;
 		default: edge_mask_reg_512p3[352] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110010011,
12'b100110100011: edge_mask_reg_512p3[353] <= 1'b1;
 		default: edge_mask_reg_512p3[353] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100101110101,
12'b100101110110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b110010000101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[354] <= 1'b1;
 		default: edge_mask_reg_512p3[354] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b110010000100,
12'b110010010100: edge_mask_reg_512p3[355] <= 1'b1;
 		default: edge_mask_reg_512p3[355] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010000111,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111010,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100101110100,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101: edge_mask_reg_512p3[356] <= 1'b1;
 		default: edge_mask_reg_512p3[356] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111101010,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101010,
12'b11011101011,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011010,
12'b11111011011,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011001010,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b100111000110,
12'b100111000111,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110110110101,
12'b110110110110,
12'b110111000110: edge_mask_reg_512p3[357] <= 1'b1;
 		default: edge_mask_reg_512p3[357] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110101,
12'b101110110,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110101,
12'b110110110,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10101110100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b10111011010,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110010,
12'b11110110011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001001,
12'b11111001010,
12'b100010010011,
12'b100010100011,
12'b100010110011: edge_mask_reg_512p3[358] <= 1'b1;
 		default: edge_mask_reg_512p3[358] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111011001,
12'b1111011010,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10111011001,
12'b10111011010,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011101001,
12'b11011101010,
12'b11111101001,
12'b11111101010,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011110111,
12'b100011111000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111110110,
12'b101111110111,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111110101,
12'b110111110110,
12'b110111110111,
12'b111011110110: edge_mask_reg_512p3[359] <= 1'b1;
 		default: edge_mask_reg_512p3[359] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110001010,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101010,
12'b100001110101,
12'b100001110110,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b101001000101,
12'b101001000110,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100100,
12'b101001100101,
12'b101001110101,
12'b101101000101,
12'b101101000110,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100100,
12'b101101100101,
12'b101101110101,
12'b110001000101,
12'b110001010101,
12'b110001100101: edge_mask_reg_512p3[360] <= 1'b1;
 		default: edge_mask_reg_512p3[360] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10100111001,
12'b10100111010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110001001,
12'b11110001010,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101101010101,
12'b101101010110,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b110001100100,
12'b110001100101,
12'b110001110100,
12'b110001110101,
12'b110101100101,
12'b110101110101: edge_mask_reg_512p3[361] <= 1'b1;
 		default: edge_mask_reg_512p3[361] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001011,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10101111101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11101011011,
12'b11101101000,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110111011,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100110,
12'b100010100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101101110110,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010100110,
12'b110101110110,
12'b110110000110,
12'b110110000111,
12'b110110010110,
12'b110110010111,
12'b111010000110: edge_mask_reg_512p3[362] <= 1'b1;
 		default: edge_mask_reg_512p3[362] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001011,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001011,
12'b1101001011,
12'b1101001100,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001011,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10101111101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110111011,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100110,
12'b100010100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010100110,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b110110000111,
12'b110110010110,
12'b110110010111,
12'b111010000111: edge_mask_reg_512p3[363] <= 1'b1;
 		default: edge_mask_reg_512p3[363] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011001,
12'b1111011010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011011000,
12'b10011011001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111011001,
12'b11001111001,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11111001001,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110000100,
12'b100110000101,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b110010010100,
12'b110010100100,
12'b110010110100: edge_mask_reg_512p3[364] <= 1'b1;
 		default: edge_mask_reg_512p3[364] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111011001,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101011000011,
12'b101011000100,
12'b101011000101,
12'b101110100100,
12'b101110100101,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010100100,
12'b110010110100: edge_mask_reg_512p3[365] <= 1'b1;
 		default: edge_mask_reg_512p3[365] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011001,
12'b11110011010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100101110011,
12'b100110000011,
12'b100110010011: edge_mask_reg_512p3[366] <= 1'b1;
 		default: edge_mask_reg_512p3[366] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011001,
12'b11110011010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100101110011,
12'b100110000011,
12'b100110010011: edge_mask_reg_512p3[367] <= 1'b1;
 		default: edge_mask_reg_512p3[367] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011001,
12'b11110011010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011: edge_mask_reg_512p3[368] <= 1'b1;
 		default: edge_mask_reg_512p3[368] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p3[369] <= 1'b1;
 		default: edge_mask_reg_512p3[369] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110011001,
12'b11110011010,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p3[370] <= 1'b1;
 		default: edge_mask_reg_512p3[370] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101001,
12'b11010101010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101101010,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110011001,
12'b11110011010,
12'b100001100011,
12'b100001110011,
12'b100001110100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100101110011,
12'b100101110100,
12'b100110000011,
12'b100110000100,
12'b101001110011,
12'b101001110100,
12'b101010000100: edge_mask_reg_512p3[371] <= 1'b1;
 		default: edge_mask_reg_512p3[371] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10101001001,
12'b10101001010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001100101,
12'b101001100110,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b101110000101,
12'b110001110100,
12'b110001110101,
12'b110010000100,
12'b110010000101: edge_mask_reg_512p3[372] <= 1'b1;
 		default: edge_mask_reg_512p3[372] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11101011001,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100,
12'b101101110100,
12'b101110000100,
12'b101110010100: edge_mask_reg_512p3[373] <= 1'b1;
 		default: edge_mask_reg_512p3[373] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001000,
12'b11011001001,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b100010000100,
12'b100010000101,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010100,
12'b110010100100: edge_mask_reg_512p3[374] <= 1'b1;
 		default: edge_mask_reg_512p3[374] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010101,
12'b1111010110,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010100,
12'b10011010101,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010100,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010011,
12'b11111010100,
12'b11111011001,
12'b11111011010,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011010011,
12'b100011010100,
12'b100110100100,
12'b100110100101,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100111000011,
12'b100111000100,
12'b100111010011,
12'b100111010100,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101110100100,
12'b101110110100: edge_mask_reg_512p3[375] <= 1'b1;
 		default: edge_mask_reg_512p3[375] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b101010100100,
12'b101010110100: edge_mask_reg_512p3[376] <= 1'b1;
 		default: edge_mask_reg_512p3[376] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110110010101,
12'b110110010110,
12'b110110100101,
12'b110110100110: edge_mask_reg_512p3[377] <= 1'b1;
 		default: edge_mask_reg_512p3[377] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110110010101,
12'b110110010110,
12'b110110100101,
12'b110110100110: edge_mask_reg_512p3[378] <= 1'b1;
 		default: edge_mask_reg_512p3[378] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011100110,
12'b110011100111,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[379] <= 1'b1;
 		default: edge_mask_reg_512p3[379] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011100110,
12'b101011100111,
12'b101011101000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011100111,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[380] <= 1'b1;
 		default: edge_mask_reg_512p3[380] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100111100111,
12'b100111101000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011100111,
12'b101011101000,
12'b101011110110,
12'b101011110111,
12'b101011111000,
12'b101111100111,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b110011100111,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111110101,
12'b110111110110,
12'b111011110110: edge_mask_reg_512p3[381] <= 1'b1;
 		default: edge_mask_reg_512p3[381] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000111,
12'b100010001000,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111110010110,
12'b111110100110: edge_mask_reg_512p3[382] <= 1'b1;
 		default: edge_mask_reg_512p3[382] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b111000000101,
12'b111000000110,
12'b111000010110: edge_mask_reg_512p3[383] <= 1'b1;
 		default: edge_mask_reg_512p3[383] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b111000000110,
12'b111000010110: edge_mask_reg_512p3[384] <= 1'b1;
 		default: edge_mask_reg_512p3[384] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b111000000110,
12'b111000010110: edge_mask_reg_512p3[385] <= 1'b1;
 		default: edge_mask_reg_512p3[385] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b111000000110,
12'b111000010110: edge_mask_reg_512p3[386] <= 1'b1;
 		default: edge_mask_reg_512p3[386] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001110100,
12'b1001110101,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000101,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101110100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11110000011,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b100010010011,
12'b100010010100,
12'b100010100011: edge_mask_reg_512p3[387] <= 1'b1;
 		default: edge_mask_reg_512p3[387] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101001001,
12'b11101001010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000101000,
12'b101000110110,
12'b101000110111,
12'b101000111000,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110110,
12'b101100110111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110000100101,
12'b110000100110,
12'b110000100111,
12'b110000110110,
12'b110000110111,
12'b110100010101,
12'b110100010110,
12'b110100100101,
12'b110100100110,
12'b110100100111,
12'b110100110101,
12'b110100110110,
12'b110100110111,
12'b111000010101,
12'b111000100101,
12'b111000100110,
12'b111000110110,
12'b111100100110,
12'b111100110110: edge_mask_reg_512p3[388] <= 1'b1;
 		default: edge_mask_reg_512p3[388] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010100,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101111000100,
12'b101111000101,
12'b101111010100,
12'b101111010101,
12'b110011010100: edge_mask_reg_512p3[389] <= 1'b1;
 		default: edge_mask_reg_512p3[389] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000111,
12'b100010001000,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000111,
12'b110101010110,
12'b110101010111,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b111001010110,
12'b111001010111,
12'b111001100110,
12'b111001110110: edge_mask_reg_512p3[390] <= 1'b1;
 		default: edge_mask_reg_512p3[390] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000111,
12'b100010001000,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000111,
12'b100110001000,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000111,
12'b101010001000,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101110000111,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001110110,
12'b110001110111,
12'b110010000111,
12'b110101010110,
12'b110101010111,
12'b110101100110,
12'b110101100111,
12'b110101110110,
12'b110101110111,
12'b111001010110,
12'b111001010111,
12'b111001100110,
12'b111001110110: edge_mask_reg_512p3[391] <= 1'b1;
 		default: edge_mask_reg_512p3[391] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111101010,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011011100,
12'b11011101010,
12'b11011101011,
12'b11110011010,
12'b11110011011,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11110111100,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111001100,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b11111011100,
12'b11111101010,
12'b11111101011,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100010111010,
12'b100010111011,
12'b100011001000,
12'b100011001001,
12'b100011001010,
12'b100011001011,
12'b100011011000,
12'b100011011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b100111000111,
12'b100111001000,
12'b100111001001,
12'b100111011000,
12'b100111011001,
12'b101010100111,
12'b101010101000,
12'b101010110111,
12'b101010111000,
12'b101010111001,
12'b101011000111,
12'b101011001000,
12'b101011001001,
12'b101011011000,
12'b101011011001,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b101110111001,
12'b101111000111,
12'b101111001000,
12'b101111001001,
12'b101111011000,
12'b101111011001,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110011000110,
12'b110011000111,
12'b110011001000,
12'b110011001001,
12'b110011010111,
12'b110011011000,
12'b110011011001,
12'b110110110110,
12'b110110110111,
12'b110110111000,
12'b110111000110,
12'b110111000111,
12'b110111001000,
12'b110111001001,
12'b110111010111,
12'b110111011000,
12'b111010110110,
12'b111010110111,
12'b111011000110,
12'b111011000111,
12'b111011001000,
12'b111011010111,
12'b111110110111,
12'b111111000111,
12'b111111001000: edge_mask_reg_512p3[392] <= 1'b1;
 		default: edge_mask_reg_512p3[392] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111000,
12'b1000111001,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000111001,
12'b10000111010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100111001,
12'b10100111010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b101000010101,
12'b101000010110,
12'b101100000110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b110000000101,
12'b110000010100,
12'b110000010101,
12'b110100000101: edge_mask_reg_512p3[393] <= 1'b1;
 		default: edge_mask_reg_512p3[393] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000101000,
12'b10000101001,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11100011001: edge_mask_reg_512p3[394] <= 1'b1;
 		default: edge_mask_reg_512p3[394] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11111011010,
12'b11111011011,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111101010,
12'b11111101011,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100111,
12'b100011101000,
12'b100011101001,
12'b100011101010,
12'b100011101011,
12'b100011110111,
12'b100011111000,
12'b100011111001,
12'b100011111010,
12'b100111010111,
12'b100111011000,
12'b100111100111,
12'b100111101000,
12'b100111101001,
12'b100111110111,
12'b100111111000,
12'b100111111001,
12'b101011011000,
12'b101011100111,
12'b101011101000,
12'b101011101001,
12'b101011110111,
12'b101011111000,
12'b101011111001,
12'b101111100110,
12'b101111100111,
12'b101111101000,
12'b101111110110,
12'b101111110111,
12'b101111111000,
12'b101111111001,
12'b110011100110,
12'b110011100111,
12'b110011101000,
12'b110011110110,
12'b110011110111,
12'b110011111000,
12'b110111100110,
12'b110111100111,
12'b110111101000,
12'b110111110110,
12'b110111110111,
12'b110111111000,
12'b111011100110,
12'b111011100111,
12'b111011101000,
12'b111011110110,
12'b111011110111,
12'b111011111000,
12'b111111100110,
12'b111111100111,
12'b111111110110,
12'b111111110111: edge_mask_reg_512p3[395] <= 1'b1;
 		default: edge_mask_reg_512p3[395] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011101001,
12'b11011101010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111011001,
12'b11111011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011010101,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000011,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010110011,
12'b101010110100,
12'b101011000011,
12'b101011000100,
12'b101011010100,
12'b101110110100,
12'b101111000100: edge_mask_reg_512p3[396] <= 1'b1;
 		default: edge_mask_reg_512p3[396] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100011000101,
12'b100011000110,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b100111000110,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000101,
12'b101011000110,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b101111000101,
12'b101111000110,
12'b110010100101,
12'b110010100110,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110110100101,
12'b110110100110,
12'b110110110101,
12'b110110110110,
12'b110111000101,
12'b110111000110: edge_mask_reg_512p3[397] <= 1'b1;
 		default: edge_mask_reg_512p3[397] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111011,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101010,
12'b10110101011,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101010,
12'b11010101011,
12'b11101011000,
12'b11101011010,
12'b11101011011,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011010,
12'b11110011011,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b101001100110,
12'b101001100111,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b110001100110,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110101100110,
12'b110101110110,
12'b110101110111,
12'b110110000110,
12'b110110000111,
12'b111010000110: edge_mask_reg_512p3[398] <= 1'b1;
 		default: edge_mask_reg_512p3[398] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100101,
12'b101100100110,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b110000100101,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100110101,
12'b110100110110,
12'b110101000101,
12'b110101000110,
12'b111000110110,
12'b111001000110: edge_mask_reg_512p3[399] <= 1'b1;
 		default: edge_mask_reg_512p3[399] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111000100,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11011000011,
12'b11011000100,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110011,
12'b11110110100,
12'b11111000011,
12'b11111000100,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100010110100,
12'b100110000011,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b101010010011,
12'b101010100011,
12'b101010110011: edge_mask_reg_512p3[400] <= 1'b1;
 		default: edge_mask_reg_512p3[400] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000110,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101110000100,
12'b101110010100,
12'b101110100100: edge_mask_reg_512p3[401] <= 1'b1;
 		default: edge_mask_reg_512p3[401] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100001000110,
12'b100001000111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b101000010101,
12'b101000010110,
12'b101000100101,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101001000110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100010101,
12'b110100100101,
12'b110100110101: edge_mask_reg_512p3[402] <= 1'b1;
 		default: edge_mask_reg_512p3[402] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100111001,
12'b11100111010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110100010101,
12'b110100100101: edge_mask_reg_512p3[403] <= 1'b1;
 		default: edge_mask_reg_512p3[403] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011010,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101011010,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101001001,
12'b11101001010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100100010100,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b101100100100,
12'b101100100101,
12'b101100100110,
12'b101100110100,
12'b101100110101,
12'b110000010100,
12'b110000010101,
12'b110000100100,
12'b110000100101,
12'b110000110100,
12'b110000110101,
12'b110100010101,
12'b110100100101: edge_mask_reg_512p3[404] <= 1'b1;
 		default: edge_mask_reg_512p3[404] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110101,
12'b100110110110,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110101,
12'b101010110110,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110101,
12'b101110110110,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110010110101,
12'b110110000100,
12'b110110010100,
12'b110110010101,
12'b110110100100,
12'b110110100101,
12'b110110110101: edge_mask_reg_512p3[405] <= 1'b1;
 		default: edge_mask_reg_512p3[405] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111010,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000010110,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100010101,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101101001,
12'b11101101010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101001000101,
12'b101001010100,
12'b101001010101,
12'b101100100100,
12'b101100110100,
12'b101101000100,
12'b101101010100: edge_mask_reg_512p3[406] <= 1'b1;
 		default: edge_mask_reg_512p3[406] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11000010110,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100010101,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101001000101,
12'b101100100100,
12'b101100110100,
12'b101101000100: edge_mask_reg_512p3[407] <= 1'b1;
 		default: edge_mask_reg_512p3[407] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101001,
12'b10101101010,
12'b11000010110,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11100010101,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010101,
12'b100001010110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101001000101,
12'b101100100100,
12'b101100110100,
12'b101100110101,
12'b101101000100,
12'b101101000101: edge_mask_reg_512p3[408] <= 1'b1;
 		default: edge_mask_reg_512p3[408] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100011000,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100010110,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010101,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000101,
12'b100001000110,
12'b100100100011,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000101,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101100100100,
12'b101100110100: edge_mask_reg_512p3[409] <= 1'b1;
 		default: edge_mask_reg_512p3[409] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101011,
12'b1100100110,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011001,
12'b11100011010,
12'b11100011011,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010100,
12'b100000010101,
12'b100000010110,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000101,
12'b100001000110,
12'b100100010100,
12'b100100100011,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101100100100,
12'b101100110100: edge_mask_reg_512p3[410] <= 1'b1;
 		default: edge_mask_reg_512p3[410] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1100100111,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100110111,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100110,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110110,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101010,
12'b10100011001,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000011001,
12'b11000011010,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11100010101,
12'b11100011001,
12'b11100011010,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101011001,
12'b11101011010,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000100,
12'b100101000101,
12'b101000100100,
12'b101000100101,
12'b101000110100,
12'b101000110101,
12'b101001000100,
12'b101100100100,
12'b101100110100: edge_mask_reg_512p3[411] <= 1'b1;
 		default: edge_mask_reg_512p3[411] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101011,
12'b10001101100,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111000,
12'b11110111010,
12'b11110111011,
12'b11111001011,
12'b100010000110,
12'b100010000111,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100010101011,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110101,
12'b101010110110,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b110010010110,
12'b110010100101,
12'b110010100110,
12'b110110100110: edge_mask_reg_512p3[412] <= 1'b1;
 		default: edge_mask_reg_512p3[412] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010101,
12'b110010110,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101110100,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110010011,
12'b100110100011: edge_mask_reg_512p3[413] <= 1'b1;
 		default: edge_mask_reg_512p3[413] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101110010,
12'b11101110011,
12'b11101111001,
12'b11101111010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b100010000011,
12'b100010010011,
12'b100010100011,
12'b100110000011,
12'b100110010011: edge_mask_reg_512p3[414] <= 1'b1;
 		default: edge_mask_reg_512p3[414] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110010,
12'b11110110011,
12'b11110111001,
12'b100010000011,
12'b100010000100,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100110010011,
12'b100110100011: edge_mask_reg_512p3[415] <= 1'b1;
 		default: edge_mask_reg_512p3[415] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101101001,
12'b10101110100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110010,
12'b11110110011,
12'b11110111001,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100110000011,
12'b100110010011,
12'b100110010100,
12'b100110100011: edge_mask_reg_512p3[416] <= 1'b1;
 		default: edge_mask_reg_512p3[416] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000110,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010110,
12'b110010111,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11110000100,
12'b11110000101,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110010,
12'b11110110011,
12'b11110111001,
12'b11110111010,
12'b100010010011,
12'b100010010100,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100110010011,
12'b100110100011: edge_mask_reg_512p3[417] <= 1'b1;
 		default: edge_mask_reg_512p3[417] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010101010,
12'b100010110011,
12'b100010110100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100: edge_mask_reg_512p3[418] <= 1'b1;
 		default: edge_mask_reg_512p3[418] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111010,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111011,
12'b1001111100,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b11000101010,
12'b11000101011,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101010,
12'b11001101011,
12'b11100101010,
12'b11100101011,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011010,
12'b11101011011,
12'b11101101011,
12'b100000110111,
12'b100000111000,
12'b100000111001,
12'b100000111010,
12'b100000111011,
12'b100001000111,
12'b100001001000,
12'b100001001001,
12'b100001001010,
12'b100001001011,
12'b100001010111,
12'b100001011000,
12'b100100101000,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010111,
12'b100101011000,
12'b101000110110,
12'b101000110111,
12'b101000111000,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001010111,
12'b101001011000,
12'b101100110110,
12'b101100110111,
12'b101100111000,
12'b101101000110,
12'b101101000111,
12'b101101001000,
12'b101101010111,
12'b110000110110,
12'b110000110111,
12'b110001000110,
12'b110001000111,
12'b110100110110,
12'b110100110111,
12'b110101000110,
12'b110101000111,
12'b111000110110,
12'b111000110111,
12'b111001000110,
12'b111001000111: edge_mask_reg_512p3[419] <= 1'b1;
 		default: edge_mask_reg_512p3[419] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011010,
12'b10110011011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101101010110,
12'b101101010111,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000111,
12'b111001100110,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111101110111: edge_mask_reg_512p3[420] <= 1'b1;
 		default: edge_mask_reg_512p3[420] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011010,
12'b10110011011,
12'b11000111010,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011010,
12'b11010011011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001010110,
12'b110001010111,
12'b110001100110,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110101010110,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000111,
12'b111001100110,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111101110111: edge_mask_reg_512p3[421] <= 1'b1;
 		default: edge_mask_reg_512p3[421] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101010,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11101011000,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011010,
12'b11110011011,
12'b100001011000,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100010001000,
12'b100010001001,
12'b100101011000,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b100110001000,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101010000111,
12'b101010001000,
12'b101101100111,
12'b101101101000,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111010000110,
12'b111010000111,
12'b111101110110,
12'b111101110111,
12'b111110000110,
12'b111110000111: edge_mask_reg_512p3[422] <= 1'b1;
 		default: edge_mask_reg_512p3[422] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10111001,
12'b110111001,
12'b110111010,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011010111,
12'b1011011000,
12'b1011011001,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11011001000,
12'b11011001001,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111100110,
12'b11111100111,
12'b11111101000,
12'b11111101001,
12'b11111110111,
12'b11111111000,
12'b11111111001,
12'b100011100110,
12'b100011100111,
12'b100011101000,
12'b100011110110,
12'b100011110111,
12'b100011111000,
12'b100111010111,
12'b100111100110,
12'b100111100111,
12'b100111101000,
12'b100111110110,
12'b100111110111,
12'b100111111000,
12'b101011010110,
12'b101011010111,
12'b101011100110,
12'b101011100111,
12'b101011110110,
12'b101011110111,
12'b101111010111,
12'b101111100101,
12'b101111100110,
12'b101111100111,
12'b101111110101,
12'b101111110110,
12'b101111110111,
12'b110011100101,
12'b110011100110,
12'b110011100111,
12'b110011110101,
12'b110011110110,
12'b110011110111,
12'b110111100101,
12'b110111100110,
12'b110111100111,
12'b110111110101,
12'b110111110110,
12'b110111110111,
12'b111011100101,
12'b111011100110,
12'b111011100111,
12'b111011110101,
12'b111011110110,
12'b111011110111,
12'b111111100101,
12'b111111100110,
12'b111111110101,
12'b111111110110: edge_mask_reg_512p3[423] <= 1'b1;
 		default: edge_mask_reg_512p3[423] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011010,
12'b11110001010,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010110111,
12'b100010111000,
12'b100010111001,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b100110110111,
12'b100110111000,
12'b100110111001,
12'b101010010111,
12'b101010011000,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101010110111,
12'b101010111000,
12'b101010111001,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b101110111001,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110010110110,
12'b110010110111,
12'b110010111000,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b110110101000,
12'b110110110110,
12'b110110110111,
12'b110110111000,
12'b111010100110,
12'b111010100111,
12'b111010101000,
12'b111010110110,
12'b111010110111,
12'b111010111000,
12'b111110100110,
12'b111110100111,
12'b111110110110,
12'b111110110111: edge_mask_reg_512p3[424] <= 1'b1;
 		default: edge_mask_reg_512p3[424] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101000,
12'b10011101001,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110101001,
12'b11110101010,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111101001,
12'b11111101010,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011010110,
12'b100011010111,
12'b100011011000,
12'b100110100111,
12'b100110110110,
12'b100110110111,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100110,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101011010101,
12'b101011010110,
12'b101011010111,
12'b101011100110,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b101111010101,
12'b101111010110,
12'b101111010111,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110011010101,
12'b110011010110,
12'b110110110101,
12'b110110110110,
12'b110111000101,
12'b110111000110,
12'b110111010101,
12'b110111010110,
12'b111010110101,
12'b111010110110,
12'b111011000101,
12'b111011000110,
12'b111011010101: edge_mask_reg_512p3[425] <= 1'b1;
 		default: edge_mask_reg_512p3[425] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101110100,
12'b10101110101,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101110100,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100110000011,
12'b100110000100,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010010011,
12'b101010010100,
12'b101010100011,
12'b101010100100: edge_mask_reg_512p3[426] <= 1'b1;
 		default: edge_mask_reg_512p3[426] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101001,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101001,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001010100,
12'b101001010101,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000011,
12'b101010000100,
12'b101101010100,
12'b101101100100,
12'b101101100101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b110001100100: edge_mask_reg_512p3[427] <= 1'b1;
 		default: edge_mask_reg_512p3[427] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b10111101001,
12'b10111101010,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011011100,
12'b11011101010,
12'b11011101011,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011010,
12'b11111011011,
12'b11111101010,
12'b11111101011,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100010111011,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100011001010,
12'b100011001011,
12'b100011010110,
12'b100011010111,
12'b100110100110,
12'b100110100111,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b100111000110,
12'b100111000111,
12'b100111001000,
12'b100111010110,
12'b100111010111,
12'b101010100110,
12'b101010100111,
12'b101010110110,
12'b101010110111,
12'b101011000110,
12'b101011000111,
12'b101011010110,
12'b101011010111,
12'b101110110110,
12'b101110110111,
12'b101111000110,
12'b101111000111,
12'b101111010110,
12'b101111010111,
12'b110010110110,
12'b110011000110,
12'b110011010110,
12'b110110110110,
12'b110111000110,
12'b110111010110: edge_mask_reg_512p3[428] <= 1'b1;
 		default: edge_mask_reg_512p3[428] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110101,
12'b100101110101,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[429] <= 1'b1;
 		default: edge_mask_reg_512p3[429] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110101,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000100,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[430] <= 1'b1;
 		default: edge_mask_reg_512p3[430] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110101,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010101010,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b101010000100,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101110010100,
12'b101110010101,
12'b101110100101: edge_mask_reg_512p3[431] <= 1'b1;
 		default: edge_mask_reg_512p3[431] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010100111,
12'b1010101000,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000110,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011010,
12'b11011011011,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111010,
12'b11110111011,
12'b11110111100,
12'b11111000110,
12'b11111001010,
12'b11111001011,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101010,
12'b100010101011,
12'b100010110101,
12'b100010110110,
12'b100010111010,
12'b100010111011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110101,
12'b101010110110,
12'b101110010101,
12'b101110100101: edge_mask_reg_512p3[432] <= 1'b1;
 		default: edge_mask_reg_512p3[432] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001101101,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011010,
12'b11010011011,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001010110,
12'b101001010111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101101111000,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110101100110,
12'b110101110110,
12'b110101110111: edge_mask_reg_512p3[433] <= 1'b1;
 		default: edge_mask_reg_512p3[433] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111000,
12'b11110111001,
12'b100010000100,
12'b100010000101,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101110010100,
12'b101110100100,
12'b101110110100,
12'b110010100100: edge_mask_reg_512p3[434] <= 1'b1;
 		default: edge_mask_reg_512p3[434] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100111,
12'b101001100110,
12'b101001100111,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110,
12'b111001110101,
12'b111001110110,
12'b111010000101,
12'b111010000110,
12'b111010010101: edge_mask_reg_512p3[435] <= 1'b1;
 		default: edge_mask_reg_512p3[435] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110010000100,
12'b110010000101,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110110000100,
12'b110110010100,
12'b110110010101: edge_mask_reg_512p3[436] <= 1'b1;
 		default: edge_mask_reg_512p3[436] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000101001,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11100011001,
12'b11100011010,
12'b101000000111,
12'b101000001000,
12'b101100000110,
12'b101100000111,
12'b110000000110,
12'b110000000111: edge_mask_reg_512p3[437] <= 1'b1;
 		default: edge_mask_reg_512p3[437] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111001,
12'b1100101001,
12'b1100101010,
12'b1100111010,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b101000000111,
12'b101000001000,
12'b101000010110,
12'b101000010111,
12'b101000011000,
12'b101100000110,
12'b101100000111,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100000111,
12'b110100010101,
12'b110100010110,
12'b111000000110,
12'b111000010110: edge_mask_reg_512p3[438] <= 1'b1;
 		default: edge_mask_reg_512p3[438] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001011,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100110,
12'b11110100111,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111010,
12'b11110111011,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100010001011,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011011,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100101110110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010010101,
12'b101010010110,
12'b101010100101,
12'b101010100110,
12'b101110000101,
12'b101110000110,
12'b101110010101,
12'b101110010110,
12'b101110100101,
12'b101110100110,
12'b110010010110: edge_mask_reg_512p3[439] <= 1'b1;
 		default: edge_mask_reg_512p3[439] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011010,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b110001010101,
12'b110001010110,
12'b110001100101,
12'b110001100110,
12'b110001110101,
12'b110101100101,
12'b110101100110: edge_mask_reg_512p3[440] <= 1'b1;
 		default: edge_mask_reg_512p3[440] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b11001111010,
12'b11001111011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11110001010,
12'b11110001011,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111010,
12'b11110111011,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010101011,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100111,
12'b100110101000,
12'b100110101001,
12'b101010010111,
12'b101010011000,
12'b101010011001,
12'b101010100111,
12'b101010101000,
12'b101010101001,
12'b101110010111,
12'b101110011000,
12'b101110011001,
12'b101110100111,
12'b101110101000,
12'b101110101001,
12'b110010010111,
12'b110010011000,
12'b110010011001,
12'b110010100111,
12'b110010101000,
12'b110010101001,
12'b110110010111,
12'b110110011000,
12'b110110100111,
12'b110110101000,
12'b110110110111,
12'b111010100111,
12'b111010101000,
12'b111010110111,
12'b111110100111,
12'b111110110111: edge_mask_reg_512p3[441] <= 1'b1;
 		default: edge_mask_reg_512p3[441] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101101110101,
12'b101101110110,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010100,
12'b101110010101,
12'b110001110101,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110110000101,
12'b110110000110: edge_mask_reg_512p3[442] <= 1'b1;
 		default: edge_mask_reg_512p3[442] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010110110,
12'b110110010110,
12'b110110010111,
12'b110110100110,
12'b110110100111,
12'b110110110110,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111010110110,
12'b111110010110,
12'b111110100110: edge_mask_reg_512p3[443] <= 1'b1;
 		default: edge_mask_reg_512p3[443] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100111,
12'b100101110110,
12'b100101110111,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100110,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110,
12'b111010000101,
12'b111010010101: edge_mask_reg_512p3[444] <= 1'b1;
 		default: edge_mask_reg_512p3[444] <= 1'b0;
 	endcase

    case({x,y,z})
12'b101001001,
12'b101001010,
12'b1000111001,
12'b1000111010,
12'b1001001010,
12'b1001001011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001010,
12'b10001001011,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001010,
12'b10101001011,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100011011,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100111010,
12'b11100111011,
12'b100000010111,
12'b100000011000,
12'b100000011001,
12'b100000011010,
12'b100000101000,
12'b100000101001,
12'b100100010111,
12'b100100011000,
12'b100100011001,
12'b100100101000,
12'b100100101001,
12'b101000000111,
12'b101000001000,
12'b101000010111,
12'b101000011000,
12'b101000011001,
12'b101000101000,
12'b101000101001,
12'b101100000111,
12'b101100001000,
12'b101100001001,
12'b101100010111,
12'b101100011000,
12'b101100011001,
12'b101100100111,
12'b101100101000,
12'b101100101001,
12'b110000000110,
12'b110000000111,
12'b110000001000,
12'b110000010111,
12'b110000011000,
12'b110000100111,
12'b110000101000,
12'b110100000110,
12'b110100000111,
12'b110100001000,
12'b110100010110,
12'b110100010111,
12'b110100011000,
12'b110100100111,
12'b110100101000,
12'b111000000110,
12'b111000000111,
12'b111000001000,
12'b111000010110,
12'b111000010111,
12'b111000011000,
12'b111100000110,
12'b111100000111,
12'b111100010111: edge_mask_reg_512p3[445] <= 1'b1;
 		default: edge_mask_reg_512p3[445] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011100110,
12'b10011100111,
12'b10011101000,
12'b10011101001,
12'b10110101001,
12'b10110101010,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010110,
12'b10111010111,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111100110,
12'b10111100111,
12'b10111101000,
12'b10111101001,
12'b10111101010,
12'b11010101001,
12'b11010101010,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010101,
12'b11011010110,
12'b11011010111,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011100101,
12'b11011100110,
12'b11011100111,
12'b11011101000,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010101,
12'b11111010110,
12'b11111010111,
12'b11111011000,
12'b11111011001,
12'b11111011010,
12'b11111100101,
12'b11111100110,
12'b11111100111,
12'b11111101001,
12'b11111101010,
12'b11111111001,
12'b100010110110,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100011010100,
12'b100011010101,
12'b100011010110,
12'b100011010111,
12'b100011100100,
12'b100011100101,
12'b100011100110,
12'b100011100111,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111000111,
12'b100111010100,
12'b100111010101,
12'b100111010110,
12'b100111010111,
12'b100111100100,
12'b100111100101,
12'b100111100110,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101011010100,
12'b101011010101,
12'b101011010110,
12'b101011100100,
12'b101011100101,
12'b101011100110,
12'b101111000100,
12'b101111000101,
12'b101111000110,
12'b101111010100,
12'b101111010101,
12'b101111010110,
12'b101111100100,
12'b101111100101,
12'b101111100110,
12'b110011000100,
12'b110011000101,
12'b110011010100,
12'b110011010101,
12'b110011100100,
12'b110011100101,
12'b110111000100,
12'b110111000101,
12'b110111010100,
12'b110111010101: edge_mask_reg_512p3[446] <= 1'b1;
 		default: edge_mask_reg_512p3[446] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11101101010,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100001110111,
12'b100001111000,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100101110111,
12'b100101111000,
12'b100110000111,
12'b100110001000,
12'b100110001001,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110011001,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010001001,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101101110111,
12'b101110000110,
12'b101110000111,
12'b101110001000,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110001110111,
12'b110010000110,
12'b110010000111,
12'b110010001000,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110000110,
12'b110110000111,
12'b110110001000,
12'b110110010110,
12'b110110010111,
12'b110110011000,
12'b110110100110,
12'b110110100111,
12'b111010000110,
12'b111010000111,
12'b111010001000,
12'b111010010110,
12'b111010010111,
12'b111010011000,
12'b111010100110,
12'b111010100111,
12'b111110000110,
12'b111110000111,
12'b111110010110,
12'b111110010111,
12'b111110100110,
12'b111110100111: edge_mask_reg_512p3[447] <= 1'b1;
 		default: edge_mask_reg_512p3[447] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001101011,
12'b10001101100,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011010,
12'b10011011011,
12'b10101101011,
12'b10101101100,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011010,
12'b10111011011,
12'b10111011100,
12'b11001101011,
12'b11001101100,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010001101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010101101,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000110,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011010,
12'b11011011011,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111010,
12'b11110111011,
12'b11110111100,
12'b11111000110,
12'b11111001010,
12'b11111001011,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011011,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101010,
12'b100010101011,
12'b100010110101,
12'b100010110110,
12'b100010111011,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b100110110101,
12'b100110110110,
12'b101010010101,
12'b101010010110,
12'b101010100101,
12'b101010100110,
12'b101010110101,
12'b101010110110,
12'b101110010101,
12'b101110010110,
12'b101110100101,
12'b101110100110,
12'b101110110110: edge_mask_reg_512p3[448] <= 1'b1;
 		default: edge_mask_reg_512p3[448] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101001010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11101011001,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110101100110,
12'b110101100111,
12'b110101110101,
12'b110101110110,
12'b110101110111,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b111001110101,
12'b111001110110,
12'b111010000101,
12'b111010000110,
12'b111010010101,
12'b111101110101,
12'b111101110110,
12'b111110000101,
12'b111110000110: edge_mask_reg_512p3[449] <= 1'b1;
 		default: edge_mask_reg_512p3[449] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111001,
12'b11010111010,
12'b11101101000,
12'b11101101001,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110,
12'b111010000101,
12'b111010010101,
12'b111010010110,
12'b111110000101: edge_mask_reg_512p3[450] <= 1'b1;
 		default: edge_mask_reg_512p3[450] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111010100,
12'b10111010101,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011010100,
12'b11011010101,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111010100,
12'b11111011001,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100110100011,
12'b100110110011,
12'b100110110100,
12'b100111000011,
12'b100111000100,
12'b101010110011,
12'b101011000011: edge_mask_reg_512p3[451] <= 1'b1;
 		default: edge_mask_reg_512p3[451] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b100111000011,
12'b101010100011,
12'b101010100100,
12'b101010110011,
12'b101010110100: edge_mask_reg_512p3[452] <= 1'b1;
 		default: edge_mask_reg_512p3[452] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000110,
12'b1011000111,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010111010,
12'b100110100011,
12'b100110100100,
12'b100110110011,
12'b100110110100,
12'b101010110100: edge_mask_reg_512p3[453] <= 1'b1;
 		default: edge_mask_reg_512p3[453] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011001,
12'b11110011010,
12'b100001010110,
12'b100001010111,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100001111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b101001010110,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b110001100101,
12'b110001100110,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111010000110: edge_mask_reg_512p3[454] <= 1'b1;
 		default: edge_mask_reg_512p3[454] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001001,
12'b11101001010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000110,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110101,
12'b101100110110,
12'b110000010101,
12'b110000010110,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110100010101,
12'b110100010110,
12'b110100100101,
12'b110100100110,
12'b110100110101,
12'b111000010110,
12'b111000100101,
12'b111000100110: edge_mask_reg_512p3[455] <= 1'b1;
 		default: edge_mask_reg_512p3[455] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010101,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010101,
12'b100000010110,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b101000010100,
12'b101000010101,
12'b101000010110,
12'b101000100101,
12'b101000100110,
12'b101100010100,
12'b101100010101,
12'b101100010110,
12'b110000000101,
12'b110000010101: edge_mask_reg_512p3[456] <= 1'b1;
 		default: edge_mask_reg_512p3[456] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010110,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100110,
12'b100100100111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100010101: edge_mask_reg_512p3[457] <= 1'b1;
 		default: edge_mask_reg_512p3[457] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010010100,
12'b11010010101,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011001,
12'b11111011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111010,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101,
12'b101110110100,
12'b101111000100: edge_mask_reg_512p3[458] <= 1'b1;
 		default: edge_mask_reg_512p3[458] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101100100,
12'b11101100101,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110101001,
12'b100001100100,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b101001110011,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[459] <= 1'b1;
 		default: edge_mask_reg_512p3[459] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b10000111011,
12'b10000111100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011010,
12'b10110011011,
12'b11001001010,
12'b11001001011,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011010,
12'b11010011011,
12'b11101001010,
12'b11101001011,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110001010,
12'b11110001011,
12'b100001011000,
12'b100001011001,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001110111,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100101010111,
12'b100101011000,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b101001010111,
12'b101001011000,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101101010111,
12'b101101011000,
12'b101101100111,
12'b101101101000,
12'b101101101001,
12'b101101110111,
12'b101101111000,
12'b101101111001,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110110000111,
12'b111001100110,
12'b111001100111,
12'b111001110110,
12'b111001110111,
12'b111101110111: edge_mask_reg_512p3[460] <= 1'b1;
 		default: edge_mask_reg_512p3[460] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011010,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110001010,
12'b10110001011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001010,
12'b11010001011,
12'b11100111010,
12'b11100111011,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101011100,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101101100,
12'b11101111010,
12'b11101111011,
12'b100001001000,
12'b100001001001,
12'b100001001010,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100101001000,
12'b100101001001,
12'b100101011000,
12'b100101011001,
12'b100101011010,
12'b100101101000,
12'b100101101001,
12'b100101101010,
12'b101001001000,
12'b101001001001,
12'b101001011000,
12'b101001011001,
12'b101001101000,
12'b101001101001,
12'b101101000111,
12'b101101001000,
12'b101101001001,
12'b101101010111,
12'b101101011000,
12'b101101011001,
12'b101101100111,
12'b101101101000,
12'b101101101001,
12'b110001000111,
12'b110001001000,
12'b110001001001,
12'b110001010111,
12'b110001011000,
12'b110001011001,
12'b110001100111,
12'b110001101000,
12'b110001101001,
12'b110101000111,
12'b110101001000,
12'b110101001001,
12'b110101010110,
12'b110101010111,
12'b110101011000,
12'b110101011001,
12'b110101100111,
12'b110101101000,
12'b110101101001,
12'b111001001000,
12'b111001010111,
12'b111001011000,
12'b111001011001,
12'b111001100111,
12'b111001101000,
12'b111001101001,
12'b111101010111,
12'b111101011000,
12'b111101100111,
12'b111101101000: edge_mask_reg_512p3[461] <= 1'b1;
 		default: edge_mask_reg_512p3[461] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001001010,
12'b11001001011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11101011010,
12'b11101011011,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011010,
12'b11110011011,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b110001100110,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110: edge_mask_reg_512p3[462] <= 1'b1;
 		default: edge_mask_reg_512p3[462] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111000,
12'b11010111001,
12'b11101101001,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101000,
12'b11110101001,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100100,
12'b100010100101,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100011,
12'b100110100100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100011,
12'b101010100100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110010000100,
12'b110010010100: edge_mask_reg_512p3[463] <= 1'b1;
 		default: edge_mask_reg_512p3[463] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111010,
12'b10110111011,
12'b11001011010,
12'b11001011011,
12'b11001100111,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111010,
12'b11010111011,
12'b11101100110,
12'b11101100111,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110101010,
12'b11110101011,
12'b100001100110,
12'b100001100111,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011010,
12'b100101100110,
12'b100101100111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b110110010110: edge_mask_reg_512p3[464] <= 1'b1;
 		default: edge_mask_reg_512p3[464] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011011000,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010010100,
12'b11010010101,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011001,
12'b11111011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101: edge_mask_reg_512p3[465] <= 1'b1;
 		default: edge_mask_reg_512p3[465] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011001,
12'b11111011010,
12'b100010100101,
12'b100010100110,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111010,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b100111010100,
12'b101010110100,
12'b101010110101,
12'b101011000100,
12'b101011000101,
12'b101110110100,
12'b101111000100: edge_mask_reg_512p3[466] <= 1'b1;
 		default: edge_mask_reg_512p3[466] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000101,
12'b110000110,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011001001,
12'b1011001010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10011001001,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b11110101010,
12'b11110110010,
12'b11110111001,
12'b100010000011,
12'b100010010011,
12'b100010100011,
12'b100110000011,
12'b100110010011: edge_mask_reg_512p3[467] <= 1'b1;
 		default: edge_mask_reg_512p3[467] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011010,
12'b10111011011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101010110101: edge_mask_reg_512p3[468] <= 1'b1;
 		default: edge_mask_reg_512p3[468] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000101100,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011010,
12'b11001011011,
12'b11100010111,
12'b11100011000,
12'b11100011010,
12'b11100011011,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101001010,
12'b11101001011,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000101001,
12'b100000101010,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100000111010,
12'b100001000110,
12'b100001000111,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000110,
12'b100101000111,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000101000,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101000111000,
12'b101100010110,
12'b101100010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b110000100101,
12'b110000100110,
12'b110000100111,
12'b110000110101,
12'b110000110110,
12'b110000110111,
12'b110100100110,
12'b110100110110,
12'b111000100110,
12'b111000110110: edge_mask_reg_512p3[469] <= 1'b1;
 		default: edge_mask_reg_512p3[469] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100101,
12'b100010100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100101,
12'b100110100110,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b110001110100,
12'b110001110101,
12'b110010000100,
12'b110010000101,
12'b110010010100: edge_mask_reg_512p3[470] <= 1'b1;
 		default: edge_mask_reg_512p3[470] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1100111011,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b10000111011,
12'b10000111100,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001101101,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101101101,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10101111101,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001011100,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11101001010,
12'b11101001011,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101101100,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110011010,
12'b11110011011,
12'b100001011000,
12'b100001011001,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100001101011,
12'b100001111000,
12'b100001111001,
12'b100001111010,
12'b100001111011,
12'b100010001000,
12'b100010001001,
12'b100010001010,
12'b100010001011,
12'b100101010111,
12'b100101011000,
12'b100101100111,
12'b100101101000,
12'b100101101001,
12'b100101110111,
12'b100101111000,
12'b100101111001,
12'b100101111010,
12'b100110001000,
12'b100110001001,
12'b101001010111,
12'b101001011000,
12'b101001100111,
12'b101001101000,
12'b101001101001,
12'b101001110111,
12'b101001111000,
12'b101001111001,
12'b101001111010,
12'b101010001000,
12'b101010001001,
12'b101101010111,
12'b101101011000,
12'b101101100111,
12'b101101101000,
12'b101101101001,
12'b101101110111,
12'b101101111000,
12'b101101111001,
12'b101110001000,
12'b101110001001,
12'b110001100111,
12'b110001101000,
12'b110001110110,
12'b110001110111,
12'b110001111000,
12'b110001111001,
12'b110010000111,
12'b110010001000,
12'b110010001001,
12'b110101100110,
12'b110101100111,
12'b110101101000,
12'b110101110110,
12'b110101110111,
12'b110101111000,
12'b110101111001,
12'b110110000111,
12'b110110001000,
12'b110110001001,
12'b111001100111,
12'b111001110111,
12'b111001111000,
12'b111010000111,
12'b111010001000,
12'b111101110111,
12'b111101111000,
12'b111110000111,
12'b111110001000: edge_mask_reg_512p3[471] <= 1'b1;
 		default: edge_mask_reg_512p3[471] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010011100,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001111010,
12'b10001111011,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111010,
12'b10101111011,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101010,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000110,
12'b11111000111,
12'b11111001000,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111011010,
12'b11111011011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100010101010,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100011000110,
12'b100011000111,
12'b100011001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b100111000110,
12'b100111000111,
12'b100111001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101011000101,
12'b101011000110,
12'b101011000111,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b101110100111,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000101,
12'b101111000110,
12'b101111000111,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110101,
12'b110010110110,
12'b110011000101,
12'b110011000110,
12'b110110100110,
12'b110110110110,
12'b110111000110: edge_mask_reg_512p3[472] <= 1'b1;
 		default: edge_mask_reg_512p3[472] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b110010000101: edge_mask_reg_512p3[473] <= 1'b1;
 		default: edge_mask_reg_512p3[473] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110110,
12'b110110111,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011010110,
12'b1011010111,
12'b1011011000,
12'b1011011001,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111010101,
12'b1111010110,
12'b1111010111,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011010100,
12'b10011010101,
12'b10011010110,
12'b10011010111,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10011101001,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111010100,
12'b10111010101,
12'b10111010110,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b10111101001,
12'b10111101010,
12'b11010010100,
12'b11010010101,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11011010100,
12'b11011010101,
12'b11011011001,
12'b11011011010,
12'b11011011011,
12'b11011101001,
12'b11011101010,
12'b11011101011,
12'b11110010101,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b11111000110,
12'b11111001001,
12'b11111001010,
12'b11111001011,
12'b11111010011,
12'b11111010100,
12'b11111010101,
12'b11111011001,
12'b11111011010,
12'b11111011011,
12'b100010100011,
12'b100010100100,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000011,
12'b100011000100,
12'b100011000101,
12'b100011001010,
12'b100011010011,
12'b100011010100,
12'b100110110011,
12'b100110110100,
12'b100111000100,
12'b100111010100: edge_mask_reg_512p3[474] <= 1'b1;
 		default: edge_mask_reg_512p3[474] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1100111001,
12'b1100111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001000100,
12'b11001000101,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11101000100,
12'b11101000101,
12'b11101001000,
12'b11101001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000100,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100,
12'b101101010100,
12'b101101100100: edge_mask_reg_512p3[475] <= 1'b1;
 		default: edge_mask_reg_512p3[475] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001000100,
12'b11001000101,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11101000100,
12'b11101001000,
12'b11101001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101000,
12'b11101101001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000100,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000100,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010011,
12'b101001100011,
12'b101001100100,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p3[476] <= 1'b1;
 		default: edge_mask_reg_512p3[476] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011001,
12'b1111011010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10011011001,
12'b10011011010,
12'b10011011011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b10111011001,
12'b10111011010,
12'b10111011011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011010,
12'b11011011011,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b11110111010,
12'b11110111011,
12'b11111001010,
12'b11111001011,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011010,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100010111010,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010100,
12'b101110010101,
12'b101110100101,
12'b101110110101: edge_mask_reg_512p3[477] <= 1'b1;
 		default: edge_mask_reg_512p3[477] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100110,
12'b1010100111,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11101111001,
12'b11101111010,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110111001,
12'b11110111010,
12'b11110111011,
12'b11111001001,
12'b11111001010,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101010100101,
12'b101010110100,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b101110100101: edge_mask_reg_512p3[478] <= 1'b1;
 		default: edge_mask_reg_512p3[478] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111000111,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000110,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011011000,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000100,
12'b100011000101,
12'b100011000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101,
12'b110110100101: edge_mask_reg_512p3[479] <= 1'b1;
 		default: edge_mask_reg_512p3[479] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001000,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1011011000,
12'b1011011001,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001000,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b1111011000,
12'b1111011001,
12'b1111011010,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011000111,
12'b10011001000,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10011011000,
12'b10011011001,
12'b10011011010,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110110110,
12'b10110110111,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111000110,
12'b10111000111,
12'b10111001000,
12'b10111001001,
12'b10111001010,
12'b10111001011,
12'b10111011000,
12'b10111011001,
12'b10111011010,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11010111000,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11011000101,
12'b11011000110,
12'b11011000111,
12'b11011001000,
12'b11011001001,
12'b11011001010,
12'b11011001011,
12'b11011011001,
12'b11011011010,
12'b11110001001,
12'b11110001010,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b11110111001,
12'b11110111010,
12'b11111000101,
12'b11111000110,
12'b11111000111,
12'b11111001001,
12'b11111001010,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100011000101,
12'b100011000110,
12'b100011000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100111000100,
12'b100111000101,
12'b100111000110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101011000100,
12'b101011000101,
12'b101011000110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110100,
12'b101110110101,
12'b101111000100,
12'b110010010100,
12'b110010010101,
12'b110010100100,
12'b110010100101,
12'b110010110100,
12'b110010110101,
12'b110110100101: edge_mask_reg_512p3[480] <= 1'b1;
 		default: edge_mask_reg_512p3[480] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001011011,
12'b10001011100,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101011011,
12'b10101011100,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10101111101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b11001011011,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11001111101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010001101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010101101,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001010,
12'b11011001011,
12'b11011001100,
12'b11101101010,
12'b11101101011,
12'b11101101100,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111010,
12'b11110111011,
12'b100001110110,
12'b100001110111,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001011,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010011011,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010101010,
12'b100010101011,
12'b100101110111,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b101110100111,
12'b110010000110,
12'b110010010110,
12'b110010100110,
12'b110110010110,
12'b110110100110: edge_mask_reg_512p3[481] <= 1'b1;
 		default: edge_mask_reg_512p3[481] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100101100101,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101010010101,
12'b101101110100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b110010010101: edge_mask_reg_512p3[482] <= 1'b1;
 		default: edge_mask_reg_512p3[482] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111001,
12'b10010111010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111001,
12'b10110111010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100101,
12'b11010101001,
12'b11010101010,
12'b11010111010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011001,
12'b11110011010,
12'b11110100101,
12'b11110101001,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100101100101,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010100,
12'b101010010101,
12'b101010100100,
12'b101101110100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101,
12'b101110100100,
12'b110010000101,
12'b110010010101: edge_mask_reg_512p3[483] <= 1'b1;
 		default: edge_mask_reg_512p3[483] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b10001001001,
12'b10001001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001100100,
12'b101001100101,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p3[484] <= 1'b1;
 		default: edge_mask_reg_512p3[484] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101001001,
12'b10101001010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100101100101,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001100101,
12'b101001100110,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110100,
12'b101101110101,
12'b101110000100,
12'b101110000101,
12'b110001110100,
12'b110001110101,
12'b110010000101: edge_mask_reg_512p3[485] <= 1'b1;
 		default: edge_mask_reg_512p3[485] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101101001,
12'b11101101010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011001,
12'b11110011010,
12'b11110101010,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010100,
12'b100010010101,
12'b100101100101,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b101001110100,
12'b101001110101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010100,
12'b101010010101,
12'b101101110100,
12'b101110000100,
12'b101110000101,
12'b101110010100,
12'b101110010101: edge_mask_reg_512p3[486] <= 1'b1;
 		default: edge_mask_reg_512p3[486] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110101001,
12'b11110101010,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101110110,
12'b100101110111,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110101,
12'b110110000101,
12'b110110000110,
12'b110110010101,
12'b110110010110,
12'b111010000101,
12'b111010000110,
12'b111010010101,
12'b111010010110,
12'b111110000110: edge_mask_reg_512p3[487] <= 1'b1;
 		default: edge_mask_reg_512p3[487] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001010,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010011010,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110110010110,
12'b110110010111,
12'b110110100110,
12'b110110100111,
12'b111010010110,
12'b111010010111,
12'b111010100110,
12'b111010100111,
12'b111110010110,
12'b111110100110: edge_mask_reg_512p3[488] <= 1'b1;
 		default: edge_mask_reg_512p3[488] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001011001,
12'b11001011010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b101001100110,
12'b101001100111,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b110001100110,
12'b110001100111,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110101110101,
12'b110101110110,
12'b110110000101,
12'b110110000110,
12'b111001110101,
12'b111001110110,
12'b111010000101,
12'b111010000110: edge_mask_reg_512p3[489] <= 1'b1;
 		default: edge_mask_reg_512p3[489] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001001,
12'b111001010,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001010,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001010,
12'b10011001011,
12'b10101101010,
12'b10101101011,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001010,
12'b10111001011,
12'b11001101010,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111001,
12'b11010111010,
12'b11010111011,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110111010,
12'b11110111011,
12'b100001110110,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b110010010101,
12'b110010100101: edge_mask_reg_512p3[490] <= 1'b1;
 		default: edge_mask_reg_512p3[490] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111011,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010101001,
12'b11010101010,
12'b11101011001,
12'b11101011010,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110011001,
12'b11110011010,
12'b100001100101,
12'b100001100110,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101100101,
12'b100101100110,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001100110,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010101,
12'b101110010110,
12'b110001110101,
12'b110001110110,
12'b110010000101,
12'b110010000110,
12'b110010010101,
12'b110010010110,
12'b110101110101,
12'b110110000101,
12'b110110000110: edge_mask_reg_512p3[491] <= 1'b1;
 		default: edge_mask_reg_512p3[491] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011000,
12'b10100011001,
12'b10100100110,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110110,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100010110,
12'b11100011001,
12'b11100011010,
12'b11100100101,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100100,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000100100,
12'b101000100101,
12'b101000100110,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100100,
12'b101100100101,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b110000100100,
12'b110000100101,
12'b110000110100,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100110101,
12'b110101000101,
12'b110101000110: edge_mask_reg_512p3[492] <= 1'b1;
 		default: edge_mask_reg_512p3[492] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1100101000,
12'b1100101001,
12'b1100101010,
12'b1100111000,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000100111,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000110111,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000011001,
12'b11000011010,
12'b11000100110,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110110,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b100000010111,
12'b100000100101,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100100101,
12'b101100100110,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b110000100101,
12'b110000100110,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100100101,
12'b110100110101,
12'b110100110110,
12'b110101000101,
12'b110101000110: edge_mask_reg_512p3[493] <= 1'b1;
 		default: edge_mask_reg_512p3[493] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b101001001,
12'b101001010,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111010,
12'b1001111011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101001100,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10000111100,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001001100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001011100,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100110111,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10100111100,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b10101001100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101011100,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110111,
12'b11000111000,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11000111100,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001001011,
12'b11001001100,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11100101001,
12'b11100101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11100111001,
12'b11100111010,
12'b11100111011,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101001010,
12'b11101001011,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101101010,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001001010,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010110,
12'b100101010111,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010110,
12'b101001010111,
12'b101100110101,
12'b101100110110,
12'b101100110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010110,
12'b101101010111,
12'b110000110101,
12'b110000110110,
12'b110001000101,
12'b110001000110,
12'b110100110101,
12'b110101000101,
12'b110101000110: edge_mask_reg_512p3[494] <= 1'b1;
 		default: edge_mask_reg_512p3[494] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011001,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011010,
12'b1001011011,
12'b1001011100,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001000,
12'b1010001010,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001011,
12'b1101011011,
12'b1101011100,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001011,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010001101,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100110,
12'b11010100111,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11101101010,
12'b11101101011,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100110,
12'b11110100111,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111011,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001010,
12'b100010001011,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011011,
12'b100010100110,
12'b100101110110,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010000110,
12'b101010010101,
12'b101010010110,
12'b101010100101,
12'b101010100110,
12'b101110000101,
12'b101110000110,
12'b101110010101,
12'b101110010110: edge_mask_reg_512p3[495] <= 1'b1;
 		default: edge_mask_reg_512p3[495] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1101001,
12'b1101010,
12'b1111001,
12'b1111010,
12'b10001001,
12'b10001010,
12'b10011010,
12'b10101001,
12'b10101010,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001000,
12'b1010001011,
12'b1010011010,
12'b1010011011,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011011,
12'b1101011100,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001011,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010001101,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010101101,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001011,
12'b11101111010,
12'b11101111011,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110100110,
12'b11110100111,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110111010,
12'b11110111011,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001011,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011011,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100101,
12'b100110100110,
12'b101010000101,
12'b101010010101,
12'b101010010110,
12'b101010100101,
12'b101010100110,
12'b101110010101,
12'b101110010110,
12'b101110100110,
12'b110010010110: edge_mask_reg_512p3[496] <= 1'b1;
 		default: edge_mask_reg_512p3[496] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100111,
12'b100100010110,
12'b100100010111,
12'b100100100110,
12'b100100100111,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100110,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100010101: edge_mask_reg_512p3[497] <= 1'b1;
 		default: edge_mask_reg_512p3[497] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100100110,
12'b100100100111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100000110,
12'b110100010101,
12'b110100010110: edge_mask_reg_512p3[498] <= 1'b1;
 		default: edge_mask_reg_512p3[498] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100010101,
12'b110100010110: edge_mask_reg_512p3[499] <= 1'b1;
 		default: edge_mask_reg_512p3[499] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100010101,
12'b110100010110: edge_mask_reg_512p3[500] <= 1'b1;
 		default: edge_mask_reg_512p3[500] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000000111,
12'b110000010101,
12'b110000010110,
12'b110000010111,
12'b110100000101,
12'b110100000110,
12'b110100010101,
12'b110100010110: edge_mask_reg_512p3[501] <= 1'b1;
 		default: edge_mask_reg_512p3[501] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b1000111001,
12'b1000111010,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100111,
12'b11100101001,
12'b11100101010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100110,
12'b100100100111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100010101: edge_mask_reg_512p3[502] <= 1'b1;
 		default: edge_mask_reg_512p3[502] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b100111001,
12'b101001001,
12'b101001010,
12'b101011010,
12'b101011011,
12'b1000111001,
12'b1000111010,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111000,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100100111,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111000,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001001,
12'b10101001010,
12'b10101001011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000110111,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11001001001,
12'b11001001010,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100100110,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100110111,
12'b11100111001,
12'b11100111010,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100000110110,
12'b100000110111,
12'b100100010101,
12'b100100010110,
12'b100100010111,
12'b100100100101,
12'b100100100110,
12'b100100100111,
12'b100100110110,
12'b100100110111,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100101,
12'b101000100110,
12'b101000100111,
12'b101000110110,
12'b101000110111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100101,
12'b101100100110,
12'b101100100111,
12'b101100110110,
12'b101100110111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110000100101,
12'b110000100110,
12'b110100000101,
12'b110100010101,
12'b110100100101: edge_mask_reg_512p3[503] <= 1'b1;
 		default: edge_mask_reg_512p3[503] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100111001,
12'b101001001,
12'b101001010,
12'b1000111001,
12'b1000111010,
12'b1001001010,
12'b1001001011,
12'b1100101001,
12'b1100101010,
12'b1100111001,
12'b1100111010,
12'b1100111011,
12'b1101001010,
12'b1101001011,
12'b10000101000,
12'b10000101001,
12'b10000101010,
12'b10000101011,
12'b10000111001,
12'b10000111010,
12'b10000111011,
12'b10001001010,
12'b10001001011,
12'b10100010111,
12'b10100011000,
12'b10100011001,
12'b10100101000,
12'b10100101001,
12'b10100101010,
12'b10100101011,
12'b10100111001,
12'b10100111010,
12'b10100111011,
12'b10101001010,
12'b10101001011,
12'b11000010111,
12'b11000011000,
12'b11000011001,
12'b11000011010,
12'b11000100111,
12'b11000101000,
12'b11000101001,
12'b11000101010,
12'b11000101011,
12'b11000111001,
12'b11000111010,
12'b11000111011,
12'b11100010110,
12'b11100010111,
12'b11100011000,
12'b11100011001,
12'b11100011010,
12'b11100011011,
12'b11100100111,
12'b11100101000,
12'b11100101001,
12'b11100101010,
12'b11100101011,
12'b11100111010,
12'b11100111011,
12'b100000010110,
12'b100000010111,
12'b100000011000,
12'b100000011010,
12'b100000100110,
12'b100000100111,
12'b100000101000,
12'b100100010110,
12'b100100010111,
12'b100100011000,
12'b100100100110,
12'b100100100111,
12'b100100101000,
12'b101000000111,
12'b101000010101,
12'b101000010110,
12'b101000010111,
12'b101000100110,
12'b101000100111,
12'b101100000110,
12'b101100000111,
12'b101100010101,
12'b101100010110,
12'b101100010111,
12'b101100100110,
12'b101100100111,
12'b110000000101,
12'b110000000110,
12'b110000010101,
12'b110000010110,
12'b110100000101,
12'b110100000110,
12'b110100010101,
12'b110100010110: edge_mask_reg_512p3[504] <= 1'b1;
 		default: edge_mask_reg_512p3[504] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101101100100,
12'b101101110100,
12'b101110000100: edge_mask_reg_512p3[505] <= 1'b1;
 		default: edge_mask_reg_512p3[505] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101000101,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101101100100,
12'b101101110100,
12'b101110000100: edge_mask_reg_512p3[506] <= 1'b1;
 		default: edge_mask_reg_512p3[506] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101000101,
12'b10101000110,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101000100,
12'b11101001001,
12'b11101001010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101011011,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101101011,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101101100100,
12'b101101110100,
12'b101110000100: edge_mask_reg_512p3[507] <= 1'b1;
 		default: edge_mask_reg_512p3[507] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b100111000,
12'b100111001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101001,
12'b110101010,
12'b110101011,
12'b1000111000,
12'b1000111001,
12'b1000111010,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001001011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1100111001,
12'b1100111010,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101001011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101010,
12'b1110101011,
12'b10000111010,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001001010,
12'b10001001011,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101001,
12'b10010101010,
12'b10101000101,
12'b10101000110,
12'b10101001000,
12'b10101001001,
12'b10101001010,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101011011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101101011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101001,
12'b10110101010,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001001000,
12'b11001001001,
12'b11001001010,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001011011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001101011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010011001,
12'b11010011010,
12'b11101000100,
12'b11101000101,
12'b11101001001,
12'b11101001010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101011001,
12'b11101011010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11101111010,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b11110001010,
12'b11110011001,
12'b11110011010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101010011,
12'b100101010100,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000100,
12'b101010000101,
12'b101101100100,
12'b101101110100,
12'b101110000100: edge_mask_reg_512p3[508] <= 1'b1;
 		default: edge_mask_reg_512p3[508] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110101,
12'b1001110110,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010111000,
12'b11010111001,
12'b11101101001,
12'b11101101010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110100011,
12'b11110100100,
12'b11110101001,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100011,
12'b100010100100,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010011,
12'b100110010100,
12'b100110100011,
12'b101001110011,
12'b101001110100,
12'b101010000011,
12'b101010000100,
12'b101010010011,
12'b101010010100: edge_mask_reg_512p3[509] <= 1'b1;
 		default: edge_mask_reg_512p3[509] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011010,
12'b1101010,
12'b1111010,
12'b10001010,
12'b10011010,
12'b10101010,
12'b101011010,
12'b101011011,
12'b101101010,
12'b101101011,
12'b101111010,
12'b101111011,
12'b110001010,
12'b110001011,
12'b110011010,
12'b110011011,
12'b110101010,
12'b110101011,
12'b110111010,
12'b110111011,
12'b111001010,
12'b1001011011,
12'b1001011100,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001011,
12'b1010001100,
12'b1010011011,
12'b1010011100,
12'b1010101010,
12'b1010101011,
12'b1010101100,
12'b1010111010,
12'b1010111011,
12'b1011001010,
12'b1011001011,
12'b1101011011,
12'b1101011100,
12'b1101101010,
12'b1101101011,
12'b1101101100,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110011100,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110101100,
12'b1110111010,
12'b1110111011,
12'b1110111100,
12'b1111001010,
12'b1111001011,
12'b10001011011,
12'b10001011100,
12'b10001101010,
12'b10001101011,
12'b10001101100,
12'b10001101101,
12'b10001111010,
12'b10001111011,
12'b10001111100,
12'b10001111101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010001100,
12'b10010001101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010011100,
12'b10010011101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010101100,
12'b10010101101,
12'b10010111010,
12'b10010111011,
12'b10010111100,
12'b10011001010,
12'b10011001011,
12'b10011001100,
12'b10101011011,
12'b10101011100,
12'b10101101010,
12'b10101101011,
12'b10101101100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10101111100,
12'b10101111101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110001100,
12'b10110001101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110011100,
12'b10110011101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110101100,
12'b10110101101,
12'b10110111010,
12'b10110111011,
12'b10110111100,
12'b10111001010,
12'b10111001011,
12'b10111001100,
12'b11001101010,
12'b11001101011,
12'b11001101100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11001111011,
12'b11001111100,
12'b11001111101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010001011,
12'b11010001100,
12'b11010001101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010011100,
12'b11010011101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010101100,
12'b11010101101,
12'b11010111010,
12'b11010111011,
12'b11010111100,
12'b11011001011,
12'b11011001100,
12'b11101101011,
12'b11101101100,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11101111010,
12'b11101111011,
12'b11101111100,
12'b11101111101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110001011,
12'b11110001100,
12'b11110001101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110011100,
12'b11110011101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101010,
12'b11110101011,
12'b11110101100,
12'b11110101101,
12'b11110111010,
12'b11110111011,
12'b11110111100,
12'b100001110111,
12'b100001111000,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010001001,
12'b100010001011,
12'b100010001100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011011,
12'b100010011100,
12'b100010100110,
12'b100010100111,
12'b100101110111,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100101,
12'b101010100110,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110100110,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111: edge_mask_reg_512p3[510] <= 1'b1;
 		default: edge_mask_reg_512p3[510] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111001000,
12'b111001001,
12'b111001010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011001001,
12'b1011001010,
12'b1011001011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1110111011,
12'b1111001001,
12'b1111001010,
12'b1111001011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010111000,
12'b10010111001,
12'b10010111010,
12'b10010111011,
12'b10011001001,
12'b10011001010,
12'b10011001011,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110011011,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110101011,
12'b10110111000,
12'b10110111001,
12'b10110111010,
12'b10110111011,
12'b10111001001,
12'b10111001010,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010011011,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010101010,
12'b11010101011,
12'b11010111001,
12'b11010111010,
12'b11011001001,
12'b11011001010,
12'b11101111001,
12'b11101111010,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110001010,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110011010,
12'b11110011011,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110101010,
12'b11110101011,
12'b11110111001,
12'b11110111010,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010011001,
12'b100010100111,
12'b100010101000,
12'b100010101001,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101110000110,
12'b101110000111,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b110010000110,
12'b110010000111,
12'b110010010110,
12'b110010010111,
12'b110010011000,
12'b110010100110,
12'b110010100111,
12'b110010101000,
12'b110110000110,
12'b110110000111,
12'b110110010101,
12'b110110010110,
12'b110110010111,
12'b110110100101,
12'b110110100110,
12'b110110100111,
12'b111010010101,
12'b111010010110,
12'b111010010111,
12'b111010100101,
12'b111010100110,
12'b111010100111,
12'b111110010110,
12'b111110100110: edge_mask_reg_512p3[511] <= 1'b1;
 		default: edge_mask_reg_512p3[511] <= 1'b0;
 	endcase

end
endmodule

