/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 5
second: 32
********************************************/

module prm_LUTX1_Ca_4_4_4_chk512p1(
	input [3:0] x,
	input [3:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p1
);

	reg [511:0] edge_mask_reg_512p1;
	assign edge_mask_512p1= edge_mask_reg_512p1;

always @( *) begin
    case({x,y,z})
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110111,
12'b100111000,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b1000110000,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110111,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101100111,
12'b1101101000,
12'b10001010111: edge_mask_reg_512p1[0] <= 1'b1;
 		default: edge_mask_reg_512p1[0] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110010,
12'b11010110011: edge_mask_reg_512p1[1] <= 1'b1;
 		default: edge_mask_reg_512p1[1] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000010,
12'b111000011,
12'b111000100,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000000,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000000,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010000111,
12'b10010001000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010111000,
12'b10010111001,
12'b10011000010,
12'b10011000011,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100: edge_mask_reg_512p1[2] <= 1'b1;
 		default: edge_mask_reg_512p1[2] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110111,
12'b10111000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110110110,
12'b110110111,
12'b110111000,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1101110111,
12'b1101111000,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100111,
12'b11010101000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100000,
12'b11110100001,
12'b11110100010: edge_mask_reg_512p1[3] <= 1'b1;
 		default: edge_mask_reg_512p1[3] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1001001: edge_mask_reg_512p1[4] <= 1'b1;
 		default: edge_mask_reg_512p1[4] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010110,
12'b110010111,
12'b110011000,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100110,
12'b1110100111,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100110,
12'b10010100111,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110100111,
12'b11001100001,
12'b11001100010,
12'b11001100110,
12'b11001100111,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11101100001,
12'b11101100010,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010111,
12'b100001100001,
12'b100001100010,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100101100001,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[5] <= 1'b1;
 		default: edge_mask_reg_512p1[5] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100000,
12'b10100001,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110000,
12'b10110001,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000000,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b111000000,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111001000,
12'b111001001,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000000,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110111,
12'b10010111000,
12'b10110100111,
12'b10110101000: edge_mask_reg_512p1[6] <= 1'b1;
 		default: edge_mask_reg_512p1[6] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b101001110011,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010010010,
12'b101010010011: edge_mask_reg_512p1[7] <= 1'b1;
 		default: edge_mask_reg_512p1[7] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10111000,
12'b10111001,
12'b10111010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1101111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110011,
12'b1110110100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010101011,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11011000010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110110001,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010110010,
12'b100010110011,
12'b100010110100,
12'b100110010100,
12'b100110010101,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110110010,
12'b100110110011,
12'b100110110100: edge_mask_reg_512p1[8] <= 1'b1;
 		default: edge_mask_reg_512p1[8] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b11010100011,
12'b11010100100,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11011000001,
12'b11011000010,
12'b11011000011,
12'b11011000100: edge_mask_reg_512p1[9] <= 1'b1;
 		default: edge_mask_reg_512p1[9] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001000011,
12'b11001000100,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101000011,
12'b11101000100,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b101001000100,
12'b101001010001,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101101010001,
12'b101101010010,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b110001010010,
12'b110001010011,
12'b110001100010,
12'b110001100011: edge_mask_reg_512p1[10] <= 1'b1;
 		default: edge_mask_reg_512p1[10] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100000,
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100100000,
12'b100100001,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b1000110000,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1100110010,
12'b1100110011,
12'b1101000010,
12'b1101000011,
12'b1101011000: edge_mask_reg_512p1[11] <= 1'b1;
 		default: edge_mask_reg_512p1[11] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110111,
12'b111000,
12'b111001,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110111,
12'b100111000,
12'b100111001,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b1000110000,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010111,
12'b1101011000,
12'b1101011001: edge_mask_reg_512p1[12] <= 1'b1;
 		default: edge_mask_reg_512p1[12] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100010,
12'b100011,
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b111000,
12'b111001,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100111000,
12'b100111001,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1100110011: edge_mask_reg_512p1[13] <= 1'b1;
 		default: edge_mask_reg_512p1[13] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b11000000,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000111,
12'b11001000,
12'b11010010,
12'b11010011,
12'b11010100,
12'b110100111,
12'b110101000,
12'b110110011,
12'b110110100,
12'b110110111,
12'b110111000,
12'b110111001,
12'b111000010,
12'b111000011,
12'b111000100: edge_mask_reg_512p1[14] <= 1'b1;
 		default: edge_mask_reg_512p1[14] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001001,
12'b1001010,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101101100,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001101100,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1101001000,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111001,
12'b10101111010,
12'b11000110110,
12'b11000110111,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001001001,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001011010,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11100110110,
12'b11100110111,
12'b11100111000,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101001001,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101011010,
12'b11101101000,
12'b11101101001,
12'b11101101010,
12'b100000110101,
12'b100000110110,
12'b100000110111,
12'b100000111000,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001001001,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001011001,
12'b100001011010,
12'b100001101000,
12'b100001101001,
12'b100001101010,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100100110111,
12'b100100111000,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101001001,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101011001,
12'b100101101000,
12'b100101101001,
12'b100101101010,
12'b101000110100,
12'b101000110101,
12'b101000110110,
12'b101000110111,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001001001,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001011001,
12'b101001101000,
12'b101001101001,
12'b101100110100,
12'b101100110101,
12'b101100110110,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101001000,
12'b101101001001,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101011001,
12'b101101101000,
12'b101101101001,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001000111,
12'b110001001000,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001011001,
12'b110001101000,
12'b110101000101,
12'b110101000110,
12'b110101000111,
12'b110101010101,
12'b110101010110,
12'b110101010111,
12'b111001010110: edge_mask_reg_512p1[15] <= 1'b1;
 		default: edge_mask_reg_512p1[15] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010101,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10111000,
12'b10111001,
12'b10111010,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110001,
12'b110110010,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110001,
12'b1010110010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110001,
12'b1110110010,
12'b1110111001,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110001,
12'b10010110010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101001,
12'b10110101010,
12'b10110110001,
12'b10110110010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11110100001,
12'b11110100010: edge_mask_reg_512p1[16] <= 1'b1;
 		default: edge_mask_reg_512p1[16] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b1001010111,
12'b1001011000,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100111,
12'b11101101000,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110111,
12'b11101111000,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011: edge_mask_reg_512p1[17] <= 1'b1;
 		default: edge_mask_reg_512p1[17] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000100,
12'b101000101,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b11001000001,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101: edge_mask_reg_512p1[18] <= 1'b1;
 		default: edge_mask_reg_512p1[18] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001: edge_mask_reg_512p1[19] <= 1'b1;
 		default: edge_mask_reg_512p1[19] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010101,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100000,
12'b10100001,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[20] <= 1'b1;
 		default: edge_mask_reg_512p1[20] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010100,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010100,
12'b11101010101,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001110010,
12'b110001110011: edge_mask_reg_512p1[21] <= 1'b1;
 		default: edge_mask_reg_512p1[21] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011001,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010101,
12'b101010010110,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010010,
12'b101110010011,
12'b101110010101,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010010,
12'b110010010011,
12'b110010010101,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110101110110,
12'b110110000010,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b110110000110: edge_mask_reg_512p1[22] <= 1'b1;
 		default: edge_mask_reg_512p1[22] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110001,
12'b10101110010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001110001,
12'b11001110010,
12'b11101010011,
12'b11101010100,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110001: edge_mask_reg_512p1[23] <= 1'b1;
 		default: edge_mask_reg_512p1[23] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110010,
12'b10110110011,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[24] <= 1'b1;
 		default: edge_mask_reg_512p1[24] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110111,
12'b1110111000,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110010,
12'b10110110011,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010110000,
12'b11010110010,
12'b11010110011,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110110000,
12'b100010010010,
12'b100010010011,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011: edge_mask_reg_512p1[25] <= 1'b1;
 		default: edge_mask_reg_512p1[25] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b1111100,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10001100,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b101111100,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110001100,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1001111100,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010001100,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1101111100,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110001100,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10101111011,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110001011,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11101110100,
12'b11101110101,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b100010000100,
12'b100010000101,
12'b100010010100,
12'b100010010101: edge_mask_reg_512p1[26] <= 1'b1;
 		default: edge_mask_reg_512p1[26] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010010,
12'b1010011,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1100001,
12'b1100010,
12'b1100011,
12'b1100100,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1110001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100000,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000111,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001110000,
12'b11001110110,
12'b11001110111,
12'b11001111000: edge_mask_reg_512p1[27] <= 1'b1;
 		default: edge_mask_reg_512p1[27] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010011,
12'b101001010100,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110011,
12'b101001110100: edge_mask_reg_512p1[28] <= 1'b1;
 		default: edge_mask_reg_512p1[28] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010010,
12'b10010011,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b110101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[29] <= 1'b1;
 		default: edge_mask_reg_512p1[29] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010010,
12'b1001010011,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010011,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[30] <= 1'b1;
 		default: edge_mask_reg_512p1[30] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100111,
12'b1010101000,
12'b1101100111,
12'b1101101000,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b10001100111,
12'b10001101000,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10101100111,
12'b10101101000,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110111,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110011000,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100101110010,
12'b100101110011,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010010,
12'b100110010011: edge_mask_reg_512p1[31] <= 1'b1;
 		default: edge_mask_reg_512p1[31] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010101,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100000,
12'b10100001,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b10111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110011,
12'b1010110100,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010: edge_mask_reg_512p1[32] <= 1'b1;
 		default: edge_mask_reg_512p1[32] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000000,
12'b10000001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11110000111,
12'b11110001000,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[33] <= 1'b1;
 		default: edge_mask_reg_512p1[33] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1001011,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100011,
12'b1100100,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1101000011,
12'b1101000100,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10001010011,
12'b10001010100,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010: edge_mask_reg_512p1[34] <= 1'b1;
 		default: edge_mask_reg_512p1[34] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010000,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100000,
12'b1100001,
12'b1100010,
12'b1100011,
12'b1100100,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100000,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10001010011,
12'b10001010100,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010: edge_mask_reg_512p1[35] <= 1'b1;
 		default: edge_mask_reg_512p1[35] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010000,
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100011,
12'b1100100,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100000,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001001000,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101101000,
12'b10101101001: edge_mask_reg_512p1[36] <= 1'b1;
 		default: edge_mask_reg_512p1[36] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b11000110001,
12'b11000110010,
12'b11001000001,
12'b11001000010,
12'b11001010001,
12'b11001010010: edge_mask_reg_512p1[37] <= 1'b1;
 		default: edge_mask_reg_512p1[37] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010101,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110001,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110000,
12'b10010110001,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010100010,
12'b11010100011,
12'b11010100100: edge_mask_reg_512p1[38] <= 1'b1;
 		default: edge_mask_reg_512p1[38] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100000,
12'b100001,
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b100100000,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b1000110010,
12'b1000110011,
12'b1001000010,
12'b1001000011,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000: edge_mask_reg_512p1[39] <= 1'b1;
 		default: edge_mask_reg_512p1[39] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10110001000,
12'b10110001001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10111000001,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110011,
12'b11010110100,
12'b11010110101: edge_mask_reg_512p1[40] <= 1'b1;
 		default: edge_mask_reg_512p1[40] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101000011,
12'b11101000100,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b100001000011,
12'b100001000100,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b101001010001,
12'b101001010010,
12'b101001010011,
12'b101001100001,
12'b101001100010: edge_mask_reg_512p1[41] <= 1'b1;
 		default: edge_mask_reg_512p1[41] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100001,
12'b10100010,
12'b10100011,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000001,
12'b110000010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100111,
12'b10110101000,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010010,
12'b11010010011,
12'b11010010111,
12'b11010011000,
12'b11010100111,
12'b11010101000: edge_mask_reg_512p1[42] <= 1'b1;
 		default: edge_mask_reg_512p1[42] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010110,
12'b1010111,
12'b1011000,
12'b1100001,
12'b1100010,
12'b1100011,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1110001,
12'b1110010,
12'b1110011,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100000,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b1001010001,
12'b1001010010,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b11001010001,
12'b11001010010,
12'b11001010111,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001110000,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11101100111: edge_mask_reg_512p1[43] <= 1'b1;
 		default: edge_mask_reg_512p1[43] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110001,
12'b10110010,
12'b10110011,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010101,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1110001001,
12'b1110001010,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111001,
12'b1110111010,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b11010100100,
12'b11010110100,
12'b11010110101: edge_mask_reg_512p1[44] <= 1'b1;
 		default: edge_mask_reg_512p1[44] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000001,
12'b10000010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010000,
12'b10010010,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100000,
12'b110100001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010111,
12'b11010011000,
12'b11010100111,
12'b11010101000,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[45] <= 1'b1;
 		default: edge_mask_reg_512p1[45] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p1[46] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010001,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100000,
12'b1100001,
12'b1100010,
12'b1100011,
12'b1100100,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101000111,
12'b101001000,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100000,
12'b101100001,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110000,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[47] <= 1'b1;
 		default: edge_mask_reg_512p1[47] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1001110111,
12'b1001111000,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010000111,
12'b11010001000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010111,
12'b11010011000,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100111,
12'b11010101000,
12'b11010110010,
12'b11010110011: edge_mask_reg_512p1[48] <= 1'b1;
 		default: edge_mask_reg_512p1[48] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010101,
12'b1010110,
12'b1010111,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1110101,
12'b1110110,
12'b1110111,
12'b10000101,
12'b10000110,
12'b10000111,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000101,
12'b110000110,
12'b110000111,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101100000,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11010000110,
12'b11010000111,
12'b11101000000,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100111,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110111,
12'b100001000001,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100101010000,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101100000,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b101001010001,
12'b101001010010,
12'b101001100000,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101101100001,
12'b101101100010,
12'b101101110001,
12'b101101110010: edge_mask_reg_512p1[49] <= 1'b1;
 		default: edge_mask_reg_512p1[49] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b100001000000,
12'b100001000001,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100101000001,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b101001010001,
12'b101001010010: edge_mask_reg_512p1[50] <= 1'b1;
 		default: edge_mask_reg_512p1[50] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1000110100,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101101001,
12'b10101101010,
12'b11000110100,
12'b11000110101,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100101000010,
12'b100101000011,
12'b100101010010,
12'b100101010011: edge_mask_reg_512p1[51] <= 1'b1;
 		default: edge_mask_reg_512p1[51] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p1[52] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010110001,
12'b11010110010,
12'b11110000011,
12'b11110000100,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110110001,
12'b11110110010,
12'b100010010011,
12'b100010100011: edge_mask_reg_512p1[53] <= 1'b1;
 		default: edge_mask_reg_512p1[53] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b101001010001,
12'b101001010010,
12'b101001100001,
12'b101001100010: edge_mask_reg_512p1[54] <= 1'b1;
 		default: edge_mask_reg_512p1[54] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100001,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010111000,
12'b10010111001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001: edge_mask_reg_512p1[55] <= 1'b1;
 		default: edge_mask_reg_512p1[55] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010110,
12'b110010111,
12'b110011000,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110111,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000111,
12'b11110001000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100101110001,
12'b100101110010,
12'b100110000001,
12'b100110000010,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[56] <= 1'b1;
 		default: edge_mask_reg_512p1[56] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001000100,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11101000011,
12'b11101000100,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010001,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101010010,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b110001100010,
12'b110001100011,
12'b110001110011: edge_mask_reg_512p1[57] <= 1'b1;
 		default: edge_mask_reg_512p1[57] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110000,
12'b10110001,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000000,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000000,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000111,
12'b111001000,
12'b111001001,
12'b1010011000,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000000,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000010,
12'b1111000011: edge_mask_reg_512p1[58] <= 1'b1;
 		default: edge_mask_reg_512p1[58] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110111,
12'b111000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b100110010,
12'b100110011,
12'b101000111,
12'b101001000,
12'b101010111,
12'b101011000: edge_mask_reg_512p1[59] <= 1'b1;
 		default: edge_mask_reg_512p1[59] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1001001,
12'b1001010,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10001000,
12'b10001001,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10000110110,
12'b10000110111,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100111,
12'b11001101000,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100100110110,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101101000011,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b110001000100,
12'b110001010100: edge_mask_reg_512p1[60] <= 1'b1;
 		default: edge_mask_reg_512p1[60] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100001,
12'b11100010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111100001,
12'b111100010,
12'b1010101000,
12'b1010101001,
12'b1010111000,
12'b1010111001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1111000011,
12'b1111000100,
12'b1111010010,
12'b1111010011,
12'b1111010100: edge_mask_reg_512p1[61] <= 1'b1;
 		default: edge_mask_reg_512p1[61] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000011,
12'b1101000100,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001011001,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b100001000011,
12'b100001000100,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b101001010001,
12'b101001010010,
12'b101001100001,
12'b101001100010: edge_mask_reg_512p1[62] <= 1'b1;
 		default: edge_mask_reg_512p1[62] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001111000,
12'b1001111001,
12'b1100110010,
12'b1100110011,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b11000110011,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11101010001: edge_mask_reg_512p1[63] <= 1'b1;
 		default: edge_mask_reg_512p1[63] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110001,
12'b11101110010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110001,
12'b100001110010,
12'b100001110100,
12'b100001110101,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001010011,
12'b101001010100,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100: edge_mask_reg_512p1[64] <= 1'b1;
 		default: edge_mask_reg_512p1[64] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100101,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10101100,
12'b10110001,
12'b10110010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b10111011,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110001,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b10010100100,
12'b10010110011,
12'b10010110100: edge_mask_reg_512p1[65] <= 1'b1;
 		default: edge_mask_reg_512p1[65] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010001000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110110010,
12'b11110110011,
12'b11110110100: edge_mask_reg_512p1[66] <= 1'b1;
 		default: edge_mask_reg_512p1[66] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000111,
12'b10110001000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010010111,
12'b11010011000,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11010110011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[67] <= 1'b1;
 		default: edge_mask_reg_512p1[67] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001111000,
12'b11001111001,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b100001010001,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001110001,
12'b100001110010: edge_mask_reg_512p1[68] <= 1'b1;
 		default: edge_mask_reg_512p1[68] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b10010101000,
12'b10010101001,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011010001,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111010001,
12'b11010110011,
12'b11010110100,
12'b11011000001,
12'b11011000010,
12'b11011000011,
12'b11011000100: edge_mask_reg_512p1[69] <= 1'b1;
 		default: edge_mask_reg_512p1[69] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110110,
12'b1110110111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10110001000,
12'b10110001001,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10110110111,
12'b10111000010,
12'b10111000011,
12'b10111000101,
12'b11010010101,
12'b11010010110,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11010110110,
12'b11010110111,
12'b11011000010,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110110001,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11111000010,
12'b11111000011,
12'b11111000100,
12'b11111000101,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010110001,
12'b100010110010,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100011000010,
12'b100011000011: edge_mask_reg_512p1[70] <= 1'b1;
 		default: edge_mask_reg_512p1[70] <= 1'b0;
 	endcase

    case({x,y,z})
12'b111000,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100010,
12'b1100011,
12'b1100100,
12'b1100101,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100010,
12'b101100011,
12'b101100100,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001: edge_mask_reg_512p1[71] <= 1'b1;
 		default: edge_mask_reg_512p1[71] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001000111,
12'b10001001000,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001001,
12'b11001000110,
12'b11001000111,
12'b11001001000,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11100110110,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b100000110101,
12'b100000110110,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100100110101,
12'b100100110110,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000011,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b110001000011,
12'b110001000100,
12'b110001000101,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101010100,
12'b110101010101,
12'b110101100100,
12'b110101100101: edge_mask_reg_512p1[72] <= 1'b1;
 		default: edge_mask_reg_512p1[72] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1000111000,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000100100,
12'b10000100101,
12'b10000100110,
12'b10000100111,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001111000,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100100111,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b11000100100,
12'b11000100101,
12'b11000100110,
12'b11000100111,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11000110111,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11100100100,
12'b11100100101,
12'b11100100110,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11100110111,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b100000100011,
12'b100000100100,
12'b100000100101,
12'b100000100110,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100100100011,
12'b100100100100,
12'b100100100101,
12'b100100110010,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b101000100011,
12'b101000100100,
12'b101000100101,
12'b101000110010,
12'b101000110011,
12'b101000110100,
12'b101000110101,
12'b101001000010,
12'b101001000011,
12'b101001000100,
12'b101100100100,
12'b101100110010,
12'b101100110011,
12'b101100110100,
12'b101100110101,
12'b101101000010,
12'b101101000011,
12'b101101000100,
12'b110000110011,
12'b110001000011: edge_mask_reg_512p1[73] <= 1'b1;
 		default: edge_mask_reg_512p1[73] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110001,
12'b1001110010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[74] <= 1'b1;
 		default: edge_mask_reg_512p1[74] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001011011,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b101001000011,
12'b101001010011,
12'b101001010100,
12'b101001100011,
12'b101101010011,
12'b101101010100: edge_mask_reg_512p1[75] <= 1'b1;
 		default: edge_mask_reg_512p1[75] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100101,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101001,
12'b11001101010,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001111001,
12'b11101010011,
12'b11101010100,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110001,
12'b11101110010: edge_mask_reg_512p1[76] <= 1'b1;
 		default: edge_mask_reg_512p1[76] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10011100,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10101100,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b10111011,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110011100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111000100,
12'b111000101,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1010111011,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110101011,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111010,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10111000010,
12'b11010100100,
12'b11010100101,
12'b11010110100,
12'b11010110101: edge_mask_reg_512p1[77] <= 1'b1;
 		default: edge_mask_reg_512p1[77] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110011,
12'b1100110100,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110011,
12'b10000110100,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b11001000001,
12'b11001000010,
12'b11001010001,
12'b11001010010: edge_mask_reg_512p1[78] <= 1'b1;
 		default: edge_mask_reg_512p1[78] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b10111011,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11010100,
12'b11010101,
12'b11010110,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110101011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b110111011,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b1010011001,
12'b1010011010,
12'b1010101001,
12'b1010101010,
12'b1010101011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011010011,
12'b10011010100: edge_mask_reg_512p1[79] <= 1'b1;
 		default: edge_mask_reg_512p1[79] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1100110101,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11100110010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100101,
12'b11101100110,
12'b100000110001,
12'b100000110010,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100001000001,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100101,
12'b100001100110,
12'b100100110010,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000001,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100010,
12'b100101100011,
12'b101000110010,
12'b101000110011,
12'b101001000001,
12'b101001000010,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001010001,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101101000010,
12'b101101000011,
12'b101101010010,
12'b101101010011: edge_mask_reg_512p1[80] <= 1'b1;
 		default: edge_mask_reg_512p1[80] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110101,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101111000,
12'b10101111001,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100110,
12'b11100110010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b100000110001,
12'b100000110010,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100001000001,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100100110010,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000001,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b101000110010,
12'b101000110011,
12'b101001000001,
12'b101001000010,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101101000010,
12'b101101000011,
12'b101101010010,
12'b101101010011: edge_mask_reg_512p1[81] <= 1'b1;
 		default: edge_mask_reg_512p1[81] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11010100,
12'b11010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111010011,
12'b111010100,
12'b111010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010000,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011100011,
12'b1011100100,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1111000000,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010000,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b1111100001,
12'b1111100010,
12'b1111100011,
12'b1111100100,
12'b10010010111,
12'b10010100111,
12'b10010101000,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000000,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011010000,
12'b10011010001,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10011010101,
12'b10011100001,
12'b10011100010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b10111000000,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111010001,
12'b10111010010,
12'b10111010011,
12'b10111010100,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11010110101,
12'b11011000001,
12'b11011000010,
12'b11011000011,
12'b11011000100,
12'b11011000101,
12'b11011010001,
12'b11011010010,
12'b11011010011,
12'b11011010100,
12'b11111000001,
12'b11111000010,
12'b11111000011,
12'b11111000100,
12'b11111010001: edge_mask_reg_512p1[82] <= 1'b1;
 		default: edge_mask_reg_512p1[82] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10100001,
12'b10100010,
12'b10100011,
12'b10100100,
12'b10100110,
12'b10100111,
12'b10101000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110110111,
12'b110111000,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010110111,
12'b1010111000,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110111,
12'b1110111000,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010100111,
12'b11010101000: edge_mask_reg_512p1[83] <= 1'b1;
 		default: edge_mask_reg_512p1[83] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101000111,
12'b101001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110001000,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101000010,
12'b11101000011,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100101010000,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101100001,
12'b100101100010,
12'b100101100011: edge_mask_reg_512p1[84] <= 1'b1;
 		default: edge_mask_reg_512p1[84] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1001011,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100100111,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111000,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101001011,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b1000010010,
12'b1000010011,
12'b1000010100,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000100110,
12'b1000100111,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1000111000,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1100010011,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100100110,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1100111000,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101011001,
12'b1101011010,
12'b10000100011,
12'b10000100100,
12'b10000100101,
12'b10000100110,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10100100011,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10101000101,
12'b10101000110,
12'b11000110101,
12'b11000110110: edge_mask_reg_512p1[85] <= 1'b1;
 		default: edge_mask_reg_512p1[85] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[86] <= 1'b1;
 		default: edge_mask_reg_512p1[86] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[87] <= 1'b1;
 		default: edge_mask_reg_512p1[87] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[88] <= 1'b1;
 		default: edge_mask_reg_512p1[88] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[89] <= 1'b1;
 		default: edge_mask_reg_512p1[89] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[90] <= 1'b1;
 		default: edge_mask_reg_512p1[90] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001101000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[91] <= 1'b1;
 		default: edge_mask_reg_512p1[91] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001101000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[92] <= 1'b1;
 		default: edge_mask_reg_512p1[92] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[93] <= 1'b1;
 		default: edge_mask_reg_512p1[93] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[94] <= 1'b1;
 		default: edge_mask_reg_512p1[94] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[95] <= 1'b1;
 		default: edge_mask_reg_512p1[95] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[96] <= 1'b1;
 		default: edge_mask_reg_512p1[96] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[97] <= 1'b1;
 		default: edge_mask_reg_512p1[97] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[98] <= 1'b1;
 		default: edge_mask_reg_512p1[98] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[99] <= 1'b1;
 		default: edge_mask_reg_512p1[99] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[100] <= 1'b1;
 		default: edge_mask_reg_512p1[100] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000010,
12'b11110000011,
12'b11110010010,
12'b11110010011: edge_mask_reg_512p1[101] <= 1'b1;
 		default: edge_mask_reg_512p1[101] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000010,
12'b11110000011,
12'b11110010010,
12'b11110010011: edge_mask_reg_512p1[102] <= 1'b1;
 		default: edge_mask_reg_512p1[102] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100100,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100010,
12'b11010100011,
12'b11110010010,
12'b11110010011: edge_mask_reg_512p1[103] <= 1'b1;
 		default: edge_mask_reg_512p1[103] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100010,
12'b11010100011,
12'b11110010010,
12'b11110010011: edge_mask_reg_512p1[104] <= 1'b1;
 		default: edge_mask_reg_512p1[104] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11110010010,
12'b11110010011: edge_mask_reg_512p1[105] <= 1'b1;
 		default: edge_mask_reg_512p1[105] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[106] <= 1'b1;
 		default: edge_mask_reg_512p1[106] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000011,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001111000,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[107] <= 1'b1;
 		default: edge_mask_reg_512p1[107] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[108] <= 1'b1;
 		default: edge_mask_reg_512p1[108] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[109] <= 1'b1;
 		default: edge_mask_reg_512p1[109] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001111000,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[110] <= 1'b1;
 		default: edge_mask_reg_512p1[110] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[111] <= 1'b1;
 		default: edge_mask_reg_512p1[111] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[112] <= 1'b1;
 		default: edge_mask_reg_512p1[112] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[113] <= 1'b1;
 		default: edge_mask_reg_512p1[113] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[114] <= 1'b1;
 		default: edge_mask_reg_512p1[114] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[115] <= 1'b1;
 		default: edge_mask_reg_512p1[115] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[116] <= 1'b1;
 		default: edge_mask_reg_512p1[116] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11101110111,
12'b11101111000,
12'b11110000010,
12'b11110000011,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[117] <= 1'b1;
 		default: edge_mask_reg_512p1[117] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[118] <= 1'b1;
 		default: edge_mask_reg_512p1[118] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[119] <= 1'b1;
 		default: edge_mask_reg_512p1[119] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[120] <= 1'b1;
 		default: edge_mask_reg_512p1[120] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[121] <= 1'b1;
 		default: edge_mask_reg_512p1[121] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[122] <= 1'b1;
 		default: edge_mask_reg_512p1[122] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[123] <= 1'b1;
 		default: edge_mask_reg_512p1[123] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[124] <= 1'b1;
 		default: edge_mask_reg_512p1[124] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[125] <= 1'b1;
 		default: edge_mask_reg_512p1[125] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[126] <= 1'b1;
 		default: edge_mask_reg_512p1[126] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[127] <= 1'b1;
 		default: edge_mask_reg_512p1[127] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[128] <= 1'b1;
 		default: edge_mask_reg_512p1[128] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[129] <= 1'b1;
 		default: edge_mask_reg_512p1[129] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[130] <= 1'b1;
 		default: edge_mask_reg_512p1[130] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[131] <= 1'b1;
 		default: edge_mask_reg_512p1[131] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[132] <= 1'b1;
 		default: edge_mask_reg_512p1[132] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[133] <= 1'b1;
 		default: edge_mask_reg_512p1[133] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[134] <= 1'b1;
 		default: edge_mask_reg_512p1[134] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[135] <= 1'b1;
 		default: edge_mask_reg_512p1[135] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[136] <= 1'b1;
 		default: edge_mask_reg_512p1[136] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[137] <= 1'b1;
 		default: edge_mask_reg_512p1[137] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[138] <= 1'b1;
 		default: edge_mask_reg_512p1[138] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[139] <= 1'b1;
 		default: edge_mask_reg_512p1[139] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[140] <= 1'b1;
 		default: edge_mask_reg_512p1[140] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[141] <= 1'b1;
 		default: edge_mask_reg_512p1[141] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[142] <= 1'b1;
 		default: edge_mask_reg_512p1[142] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[143] <= 1'b1;
 		default: edge_mask_reg_512p1[143] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[144] <= 1'b1;
 		default: edge_mask_reg_512p1[144] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[145] <= 1'b1;
 		default: edge_mask_reg_512p1[145] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[146] <= 1'b1;
 		default: edge_mask_reg_512p1[146] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[147] <= 1'b1;
 		default: edge_mask_reg_512p1[147] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[148] <= 1'b1;
 		default: edge_mask_reg_512p1[148] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[149] <= 1'b1;
 		default: edge_mask_reg_512p1[149] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[150] <= 1'b1;
 		default: edge_mask_reg_512p1[150] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[151] <= 1'b1;
 		default: edge_mask_reg_512p1[151] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[152] <= 1'b1;
 		default: edge_mask_reg_512p1[152] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[153] <= 1'b1;
 		default: edge_mask_reg_512p1[153] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110011000,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[154] <= 1'b1;
 		default: edge_mask_reg_512p1[154] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[155] <= 1'b1;
 		default: edge_mask_reg_512p1[155] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000: edge_mask_reg_512p1[156] <= 1'b1;
 		default: edge_mask_reg_512p1[156] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000: edge_mask_reg_512p1[157] <= 1'b1;
 		default: edge_mask_reg_512p1[157] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b11001101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000: edge_mask_reg_512p1[158] <= 1'b1;
 		default: edge_mask_reg_512p1[158] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[159] <= 1'b1;
 		default: edge_mask_reg_512p1[159] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[160] <= 1'b1;
 		default: edge_mask_reg_512p1[160] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101011000,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[161] <= 1'b1;
 		default: edge_mask_reg_512p1[161] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101011000,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001011000,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[162] <= 1'b1;
 		default: edge_mask_reg_512p1[162] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[163] <= 1'b1;
 		default: edge_mask_reg_512p1[163] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[164] <= 1'b1;
 		default: edge_mask_reg_512p1[164] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100010,
12'b11001100011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[165] <= 1'b1;
 		default: edge_mask_reg_512p1[165] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100010,
12'b11001100011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101111000: edge_mask_reg_512p1[166] <= 1'b1;
 		default: edge_mask_reg_512p1[166] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100010,
12'b11001100011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001: edge_mask_reg_512p1[167] <= 1'b1;
 		default: edge_mask_reg_512p1[167] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010001000: edge_mask_reg_512p1[168] <= 1'b1;
 		default: edge_mask_reg_512p1[168] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[169] <= 1'b1;
 		default: edge_mask_reg_512p1[169] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[170] <= 1'b1;
 		default: edge_mask_reg_512p1[170] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001010010,
12'b11001010011,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[171] <= 1'b1;
 		default: edge_mask_reg_512p1[171] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010100,
12'b1001010101,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001010010,
12'b11001010011,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101110010,
12'b11101110011: edge_mask_reg_512p1[172] <= 1'b1;
 		default: edge_mask_reg_512p1[172] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010100,
12'b1001010101,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110001000,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011,
12'b11101110010,
12'b11101110011: edge_mask_reg_512p1[173] <= 1'b1;
 		default: edge_mask_reg_512p1[173] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011,
12'b11101110010,
12'b11101110011: edge_mask_reg_512p1[174] <= 1'b1;
 		default: edge_mask_reg_512p1[174] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011,
12'b11101110010,
12'b11101110011: edge_mask_reg_512p1[175] <= 1'b1;
 		default: edge_mask_reg_512p1[175] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[176] <= 1'b1;
 		default: edge_mask_reg_512p1[176] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010010,
12'b11101010011,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[177] <= 1'b1;
 		default: edge_mask_reg_512p1[177] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010010,
12'b11101010011,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[178] <= 1'b1;
 		default: edge_mask_reg_512p1[178] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000010,
12'b10001000011,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101010010,
12'b11101010011,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[179] <= 1'b1;
 		default: edge_mask_reg_512p1[179] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10001000,
12'b101001000,
12'b101001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000100,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11101010010,
12'b11101010011,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[180] <= 1'b1;
 		default: edge_mask_reg_512p1[180] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101001000,
12'b101001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[181] <= 1'b1;
 		default: edge_mask_reg_512p1[181] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[182] <= 1'b1;
 		default: edge_mask_reg_512p1[182] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110010,
12'b11101110011,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[183] <= 1'b1;
 		default: edge_mask_reg_512p1[183] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[184] <= 1'b1;
 		default: edge_mask_reg_512p1[184] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[185] <= 1'b1;
 		default: edge_mask_reg_512p1[185] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[186] <= 1'b1;
 		default: edge_mask_reg_512p1[186] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[187] <= 1'b1;
 		default: edge_mask_reg_512p1[187] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[188] <= 1'b1;
 		default: edge_mask_reg_512p1[188] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010011000,
12'b11010011001,
12'b11110000000,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[189] <= 1'b1;
 		default: edge_mask_reg_512p1[189] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11110000000,
12'b11110000001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[190] <= 1'b1;
 		default: edge_mask_reg_512p1[190] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010011000,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b100010000000,
12'b100010000001: edge_mask_reg_512p1[191] <= 1'b1;
 		default: edge_mask_reg_512p1[191] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101110010,
12'b1101110011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001101000,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010010001: edge_mask_reg_512p1[192] <= 1'b1;
 		default: edge_mask_reg_512p1[192] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001101000,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b100001110010,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100110010001: edge_mask_reg_512p1[193] <= 1'b1;
 		default: edge_mask_reg_512p1[193] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100110000001,
12'b100110010001: edge_mask_reg_512p1[194] <= 1'b1;
 		default: edge_mask_reg_512p1[194] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100110000001,
12'b100110000011,
12'b100110000100,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[195] <= 1'b1;
 		default: edge_mask_reg_512p1[195] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010001,
12'b100110010010,
12'b100110010011: edge_mask_reg_512p1[196] <= 1'b1;
 		default: edge_mask_reg_512p1[196] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b101010010001,
12'b101010010010: edge_mask_reg_512p1[197] <= 1'b1;
 		default: edge_mask_reg_512p1[197] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100010,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100001,
12'b100110100010,
12'b101010000011,
12'b101010000100,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010100010: edge_mask_reg_512p1[198] <= 1'b1;
 		default: edge_mask_reg_512p1[198] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100010,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100001,
12'b100110100010,
12'b101010000011,
12'b101010000100,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010100010: edge_mask_reg_512p1[199] <= 1'b1;
 		default: edge_mask_reg_512p1[199] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100010,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100010,
12'b101010100011,
12'b101110010001: edge_mask_reg_512p1[200] <= 1'b1;
 		default: edge_mask_reg_512p1[200] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100010,
12'b101010100011,
12'b101110010001,
12'b101110010010,
12'b101110010100,
12'b101110100010: edge_mask_reg_512p1[201] <= 1'b1;
 		default: edge_mask_reg_512p1[201] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010: edge_mask_reg_512p1[202] <= 1'b1;
 		default: edge_mask_reg_512p1[202] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b101110100100: edge_mask_reg_512p1[203] <= 1'b1;
 		default: edge_mask_reg_512p1[203] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b110010100010: edge_mask_reg_512p1[204] <= 1'b1;
 		default: edge_mask_reg_512p1[204] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b110010100010,
12'b110010100011: edge_mask_reg_512p1[205] <= 1'b1;
 		default: edge_mask_reg_512p1[205] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110011,
12'b110010100010,
12'b110010100011: edge_mask_reg_512p1[206] <= 1'b1;
 		default: edge_mask_reg_512p1[206] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110011,
12'b110010100010,
12'b110010100011,
12'b110010100100: edge_mask_reg_512p1[207] <= 1'b1;
 		default: edge_mask_reg_512p1[207] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110011,
12'b101110110100,
12'b110010100011,
12'b110010100100: edge_mask_reg_512p1[208] <= 1'b1;
 		default: edge_mask_reg_512p1[208] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000101,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b101010000100,
12'b101010000101,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110011,
12'b101110110100,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011: edge_mask_reg_512p1[209] <= 1'b1;
 		default: edge_mask_reg_512p1[209] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000110,
12'b11110000111,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010000110,
12'b100010000111,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011,
12'b110010110100: edge_mask_reg_512p1[210] <= 1'b1;
 		default: edge_mask_reg_512p1[210] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111001,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000111,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010000110,
12'b100010000111,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100110000110,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011,
12'b110010110100,
12'b110110110100: edge_mask_reg_512p1[211] <= 1'b1;
 		default: edge_mask_reg_512p1[211] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110011,
12'b110010110100,
12'b110010110101,
12'b110110100100,
12'b110110110100: edge_mask_reg_512p1[212] <= 1'b1;
 		default: edge_mask_reg_512p1[212] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p1[213] <= 1'b1;
 		default: edge_mask_reg_512p1[213] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p1[214] <= 1'b1;
 		default: edge_mask_reg_512p1[214] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110111,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b110010010110,
12'b110010010111,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b110110110110: edge_mask_reg_512p1[215] <= 1'b1;
 		default: edge_mask_reg_512p1[215] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010001,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100010,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110011,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b110110110110: edge_mask_reg_512p1[216] <= 1'b1;
 		default: edge_mask_reg_512p1[216] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111001,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110010,
12'b11110110011,
12'b11110110100,
12'b11110110101,
12'b11110110110,
12'b11110110111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110000,
12'b100010110001,
12'b100010110010,
12'b100010110011,
12'b100010110100,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100000,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110000,
12'b100110110001,
12'b100110110010,
12'b100110110011,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100000,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110000,
12'b101010110001,
12'b101010110010,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110011000,
12'b101110100000,
12'b101110100001,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110101000,
12'b101110110000,
12'b101110110001,
12'b101110110010,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101110111000,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100001,
12'b110010100010,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110001,
12'b110010110010,
12'b110010110011,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110110100011,
12'b110110100100,
12'b110110100101,
12'b110110110011,
12'b110110110100,
12'b110110110101,
12'b110110110110: edge_mask_reg_512p1[217] <= 1'b1;
 		default: edge_mask_reg_512p1[217] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[218] <= 1'b1;
 		default: edge_mask_reg_512p1[218] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[219] <= 1'b1;
 		default: edge_mask_reg_512p1[219] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[220] <= 1'b1;
 		default: edge_mask_reg_512p1[220] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[221] <= 1'b1;
 		default: edge_mask_reg_512p1[221] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[222] <= 1'b1;
 		default: edge_mask_reg_512p1[222] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[223] <= 1'b1;
 		default: edge_mask_reg_512p1[223] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11101111001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[224] <= 1'b1;
 		default: edge_mask_reg_512p1[224] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11101111001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[225] <= 1'b1;
 		default: edge_mask_reg_512p1[225] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11101111001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[226] <= 1'b1;
 		default: edge_mask_reg_512p1[226] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101111000,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[227] <= 1'b1;
 		default: edge_mask_reg_512p1[227] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[228] <= 1'b1;
 		default: edge_mask_reg_512p1[228] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[229] <= 1'b1;
 		default: edge_mask_reg_512p1[229] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000: edge_mask_reg_512p1[230] <= 1'b1;
 		default: edge_mask_reg_512p1[230] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011: edge_mask_reg_512p1[231] <= 1'b1;
 		default: edge_mask_reg_512p1[231] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100: edge_mask_reg_512p1[232] <= 1'b1;
 		default: edge_mask_reg_512p1[232] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100: edge_mask_reg_512p1[233] <= 1'b1;
 		default: edge_mask_reg_512p1[233] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100101110000,
12'b100101110001,
12'b100101110011,
12'b100110000000,
12'b100110000001,
12'b100110000011: edge_mask_reg_512p1[234] <= 1'b1;
 		default: edge_mask_reg_512p1[234] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[235] <= 1'b1;
 		default: edge_mask_reg_512p1[235] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[236] <= 1'b1;
 		default: edge_mask_reg_512p1[236] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b101001110001,
12'b101010000001: edge_mask_reg_512p1[237] <= 1'b1;
 		default: edge_mask_reg_512p1[237] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p1[238] <= 1'b1;
 		default: edge_mask_reg_512p1[238] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p1[239] <= 1'b1;
 		default: edge_mask_reg_512p1[239] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p1[240] <= 1'b1;
 		default: edge_mask_reg_512p1[240] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110001,
12'b101101110010,
12'b101110000001,
12'b101110000010: edge_mask_reg_512p1[241] <= 1'b1;
 		default: edge_mask_reg_512p1[241] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100: edge_mask_reg_512p1[242] <= 1'b1;
 		default: edge_mask_reg_512p1[242] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100: edge_mask_reg_512p1[243] <= 1'b1;
 		default: edge_mask_reg_512p1[243] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101: edge_mask_reg_512p1[244] <= 1'b1;
 		default: edge_mask_reg_512p1[244] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110010,
12'b110010000010: edge_mask_reg_512p1[245] <= 1'b1;
 		default: edge_mask_reg_512p1[245] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110010,
12'b110001110011,
12'b110010000010,
12'b110010000011: edge_mask_reg_512p1[246] <= 1'b1;
 		default: edge_mask_reg_512p1[246] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101001,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101: edge_mask_reg_512p1[247] <= 1'b1;
 		default: edge_mask_reg_512p1[247] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101: edge_mask_reg_512p1[248] <= 1'b1;
 		default: edge_mask_reg_512p1[248] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101: edge_mask_reg_512p1[249] <= 1'b1;
 		default: edge_mask_reg_512p1[249] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001110000,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000000,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110000,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000000,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b110001110001,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000001,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101: edge_mask_reg_512p1[250] <= 1'b1;
 		default: edge_mask_reg_512p1[250] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[251] <= 1'b1;
 		default: edge_mask_reg_512p1[251] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[252] <= 1'b1;
 		default: edge_mask_reg_512p1[252] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[253] <= 1'b1;
 		default: edge_mask_reg_512p1[253] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[254] <= 1'b1;
 		default: edge_mask_reg_512p1[254] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110000,
12'b11101110001,
12'b11101111000,
12'b11101111001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[255] <= 1'b1;
 		default: edge_mask_reg_512p1[255] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110000,
12'b11101110001,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[256] <= 1'b1;
 		default: edge_mask_reg_512p1[256] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b100001110000,
12'b100001110001: edge_mask_reg_512p1[257] <= 1'b1;
 		default: edge_mask_reg_512p1[257] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110100,
12'b1001110101,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100010000000,
12'b100010000001: edge_mask_reg_512p1[258] <= 1'b1;
 		default: edge_mask_reg_512p1[258] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110101,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100101110001: edge_mask_reg_512p1[259] <= 1'b1;
 		default: edge_mask_reg_512p1[259] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000001,
12'b100010000010,
12'b100101110001,
12'b100101110010,
12'b100110000001: edge_mask_reg_512p1[260] <= 1'b1;
 		default: edge_mask_reg_512p1[260] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000001,
12'b100010000010,
12'b100101100011,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100110000001,
12'b101001110001: edge_mask_reg_512p1[261] <= 1'b1;
 		default: edge_mask_reg_512p1[261] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000001,
12'b100010000010,
12'b100101100011,
12'b100101100100,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b101001110001,
12'b101001110010,
12'b101010000001: edge_mask_reg_512p1[262] <= 1'b1;
 		default: edge_mask_reg_512p1[262] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b101001110001,
12'b101001110010,
12'b101010000001: edge_mask_reg_512p1[263] <= 1'b1;
 		default: edge_mask_reg_512p1[263] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11110000010,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001: edge_mask_reg_512p1[264] <= 1'b1;
 		default: edge_mask_reg_512p1[264] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101101110001,
12'b101101110010: edge_mask_reg_512p1[265] <= 1'b1;
 		default: edge_mask_reg_512p1[265] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100010,
12'b101101110001,
12'b101101110010: edge_mask_reg_512p1[266] <= 1'b1;
 		default: edge_mask_reg_512p1[266] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b110001110010: edge_mask_reg_512p1[267] <= 1'b1;
 		default: edge_mask_reg_512p1[267] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b110001100010,
12'b110001110010: edge_mask_reg_512p1[268] <= 1'b1;
 		default: edge_mask_reg_512p1[268] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010001000,
12'b11010001001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010100,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001110010,
12'b110001110011: edge_mask_reg_512p1[269] <= 1'b1;
 		default: edge_mask_reg_512p1[269] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001110010,
12'b110001110011: edge_mask_reg_512p1[270] <= 1'b1;
 		default: edge_mask_reg_512p1[270] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010100,
12'b101101010101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110101100011: edge_mask_reg_512p1[271] <= 1'b1;
 		default: edge_mask_reg_512p1[271] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010100,
12'b101101010101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110101100011: edge_mask_reg_512p1[272] <= 1'b1;
 		default: edge_mask_reg_512p1[272] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[273] <= 1'b1;
 		default: edge_mask_reg_512p1[273] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110100,
12'b101001110110,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110011,
12'b101101110100,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[274] <= 1'b1;
 		default: edge_mask_reg_512p1[274] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110011,
12'b101101110100,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101010011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[275] <= 1'b1;
 		default: edge_mask_reg_512p1[275] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110111,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101000101,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b101001000101,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101010011,
12'b110101010100,
12'b110101100011,
12'b110101100100,
12'b110101100101: edge_mask_reg_512p1[276] <= 1'b1;
 		default: edge_mask_reg_512p1[276] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110111,
12'b100001000110,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110111,
12'b100101000101,
12'b100101000110,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101100011,
12'b110101100100,
12'b110101100101: edge_mask_reg_512p1[277] <= 1'b1;
 		default: edge_mask_reg_512p1[277] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001001,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110111,
12'b100001000110,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000101,
12'b101101000110,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101100011,
12'b110101100100,
12'b110101100101: edge_mask_reg_512p1[278] <= 1'b1;
 		default: edge_mask_reg_512p1[278] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001001,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101010100,
12'b110101010101,
12'b110101100100,
12'b110101100101: edge_mask_reg_512p1[279] <= 1'b1;
 		default: edge_mask_reg_512p1[279] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001000111,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101000100,
12'b110101000101,
12'b110101010100,
12'b110101010101,
12'b110101100100: edge_mask_reg_512p1[280] <= 1'b1;
 		default: edge_mask_reg_512p1[280] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11101000111,
12'b11101001000,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001000111,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100110,
12'b110001100111,
12'b110101000100,
12'b110101000101,
12'b110101000110,
12'b110101010100,
12'b110101010101,
12'b110101010110: edge_mask_reg_512p1[281] <= 1'b1;
 		default: edge_mask_reg_512p1[281] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101000111,
12'b11101001000,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000001,
12'b100110000010,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000001,
12'b101010000010,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000010,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001000111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110101000100,
12'b110101000101,
12'b110101000110,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101010110,
12'b110101100011,
12'b110101100100,
12'b110101100101,
12'b110101110010,
12'b110101110011: edge_mask_reg_512p1[282] <= 1'b1;
 		default: edge_mask_reg_512p1[282] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001001,
12'b1010001010,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101001000,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101011001,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001000111,
12'b100001001000,
12'b100001010000,
12'b100001010001,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001101001,
12'b100101000000,
12'b100101000001,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101001000,
12'b100101010000,
12'b100101010001,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b101001000000,
12'b101001000001,
12'b101001000010,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001001000,
12'b101001010000,
12'b101001010001,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101101000000,
12'b101101000001,
12'b101101000010,
12'b101101000011,
12'b101101000100,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010000,
12'b101101010001,
12'b101101010010,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101011000,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101101000,
12'b110001000001,
12'b110001000010,
12'b110001000011,
12'b110001000100,
12'b110001000101,
12'b110001000110,
12'b110001000111,
12'b110001010001,
12'b110001010010,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001011000,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110101000011,
12'b110101000100,
12'b110101000101,
12'b110101000110,
12'b110101010010,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101010110: edge_mask_reg_512p1[283] <= 1'b1;
 		default: edge_mask_reg_512p1[283] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[284] <= 1'b1;
 		default: edge_mask_reg_512p1[284] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[285] <= 1'b1;
 		default: edge_mask_reg_512p1[285] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001101000,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[286] <= 1'b1;
 		default: edge_mask_reg_512p1[286] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[287] <= 1'b1;
 		default: edge_mask_reg_512p1[287] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[288] <= 1'b1;
 		default: edge_mask_reg_512p1[288] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[289] <= 1'b1;
 		default: edge_mask_reg_512p1[289] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100010,
12'b10010100011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[290] <= 1'b1;
 		default: edge_mask_reg_512p1[290] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001: edge_mask_reg_512p1[291] <= 1'b1;
 		default: edge_mask_reg_512p1[291] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010101000: edge_mask_reg_512p1[292] <= 1'b1;
 		default: edge_mask_reg_512p1[292] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010101000: edge_mask_reg_512p1[293] <= 1'b1;
 		default: edge_mask_reg_512p1[293] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010101000: edge_mask_reg_512p1[294] <= 1'b1;
 		default: edge_mask_reg_512p1[294] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000100,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110111000,
12'b1110111001,
12'b10010000010,
12'b10010000011,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011: edge_mask_reg_512p1[295] <= 1'b1;
 		default: edge_mask_reg_512p1[295] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100: edge_mask_reg_512p1[296] <= 1'b1;
 		default: edge_mask_reg_512p1[296] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101: edge_mask_reg_512p1[297] <= 1'b1;
 		default: edge_mask_reg_512p1[297] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010001000,
12'b10010001001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010111000,
12'b10010111001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110000,
12'b11010110001,
12'b11010110011: edge_mask_reg_512p1[298] <= 1'b1;
 		default: edge_mask_reg_512p1[298] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011: edge_mask_reg_512p1[299] <= 1'b1;
 		default: edge_mask_reg_512p1[299] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110101,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10011000000,
12'b10011000001,
12'b10011000011,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100: edge_mask_reg_512p1[300] <= 1'b1;
 		default: edge_mask_reg_512p1[300] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000010,
12'b111000011,
12'b111000100,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000000,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10011000000,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10110011000,
12'b10110011001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100: edge_mask_reg_512p1[301] <= 1'b1;
 		default: edge_mask_reg_512p1[301] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000000,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b11010110011,
12'b11010110100: edge_mask_reg_512p1[302] <= 1'b1;
 		default: edge_mask_reg_512p1[302] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010011000,
12'b10010011001,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10110100011,
12'b10110100100,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b11010110011: edge_mask_reg_512p1[303] <= 1'b1;
 		default: edge_mask_reg_512p1[303] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111010011,
12'b111010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010011,
12'b1011010100,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b10010101000,
12'b10010101001,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10110110011,
12'b10110110100,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100: edge_mask_reg_512p1[304] <= 1'b1;
 		default: edge_mask_reg_512p1[304] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110011,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11010011,
12'b11010100,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111010011,
12'b111010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1110011000,
12'b1110011001,
12'b1110100100,
12'b1110100101,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10110110011,
12'b10110110100,
12'b10111000001,
12'b10111000011,
12'b10111000100: edge_mask_reg_512p1[305] <= 1'b1;
 		default: edge_mask_reg_512p1[305] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001001,
12'b11010011,
12'b11010100,
12'b11010101,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011010001,
12'b10011010010,
12'b10111000011,
12'b10111000100: edge_mask_reg_512p1[306] <= 1'b1;
 		default: edge_mask_reg_512p1[306] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b1010011000,
12'b1010011001,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1110101000,
12'b1110101001,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011010001,
12'b10011010010: edge_mask_reg_512p1[307] <= 1'b1;
 		default: edge_mask_reg_512p1[307] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1110110100,
12'b1110110101,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b10011000011,
12'b10011000100,
12'b10011010100: edge_mask_reg_512p1[308] <= 1'b1;
 		default: edge_mask_reg_512p1[308] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100001,
12'b11100010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111100001,
12'b111100010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b10011000011,
12'b10011000100: edge_mask_reg_512p1[309] <= 1'b1;
 		default: edge_mask_reg_512p1[309] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100001,
12'b11100010,
12'b11100011,
12'b11100100,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100001,
12'b111100010,
12'b111100011,
12'b1010101000,
12'b1010101001,
12'b1010111000,
12'b1010111001,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111010011,
12'b1111010100,
12'b1111010101: edge_mask_reg_512p1[310] <= 1'b1;
 		default: edge_mask_reg_512p1[310] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100010,
12'b11100011,
12'b11100100,
12'b11100101,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100010,
12'b111100011,
12'b111100100,
12'b111100101,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011100010,
12'b1111010100: edge_mask_reg_512p1[311] <= 1'b1;
 		default: edge_mask_reg_512p1[311] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100010,
12'b11100011,
12'b11100100,
12'b11100101,
12'b110101000,
12'b110101001,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100010,
12'b111100011,
12'b111100100,
12'b111100101,
12'b1011000101,
12'b1011010011,
12'b1011010100,
12'b1011010101: edge_mask_reg_512p1[312] <= 1'b1;
 		default: edge_mask_reg_512p1[312] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11010111,
12'b11100010,
12'b11100011,
12'b11100100,
12'b11100101,
12'b110101000,
12'b110101001,
12'b110111000,
12'b110111001,
12'b111000101,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100010,
12'b111100011,
12'b111100100,
12'b111100101: edge_mask_reg_512p1[313] <= 1'b1;
 		default: edge_mask_reg_512p1[313] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11010111,
12'b11100010,
12'b11100011,
12'b11100100,
12'b11100101,
12'b111010100,
12'b111010101,
12'b111100100,
12'b111100101: edge_mask_reg_512p1[314] <= 1'b1;
 		default: edge_mask_reg_512p1[314] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11010111,
12'b11100001,
12'b11100010,
12'b11100011,
12'b11100100,
12'b11100101,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100001,
12'b111100010,
12'b111100011,
12'b111100100,
12'b111100101,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1011100010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1110111010,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10010111001,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011010001,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10111000001,
12'b10111000010,
12'b10111000011,
12'b10111000100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[315] <= 1'b1;
 		default: edge_mask_reg_512p1[315] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10101000,
12'b10101001,
12'b10110111,
12'b10111000,
12'b10111001,
12'b11001000,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100011,
12'b11100100,
12'b11100101: edge_mask_reg_512p1[316] <= 1'b1;
 		default: edge_mask_reg_512p1[316] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[317] <= 1'b1;
 		default: edge_mask_reg_512p1[317] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11110000111,
12'b11110001000: edge_mask_reg_512p1[318] <= 1'b1;
 		default: edge_mask_reg_512p1[318] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000: edge_mask_reg_512p1[319] <= 1'b1;
 		default: edge_mask_reg_512p1[319] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101011000,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[320] <= 1'b1;
 		default: edge_mask_reg_512p1[320] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101110111,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[321] <= 1'b1;
 		default: edge_mask_reg_512p1[321] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101111000,
12'b11101111001: edge_mask_reg_512p1[322] <= 1'b1;
 		default: edge_mask_reg_512p1[322] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001: edge_mask_reg_512p1[323] <= 1'b1;
 		default: edge_mask_reg_512p1[323] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010010,
12'b1001010011,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010010,
12'b10101010011,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100010,
12'b11001100011,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[324] <= 1'b1;
 		default: edge_mask_reg_512p1[324] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[325] <= 1'b1;
 		default: edge_mask_reg_512p1[325] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010001000,
12'b1010001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[326] <= 1'b1;
 		default: edge_mask_reg_512p1[326] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[327] <= 1'b1;
 		default: edge_mask_reg_512p1[327] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b101001000,
12'b101001001,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000010,
12'b10001000011,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001: edge_mask_reg_512p1[328] <= 1'b1;
 		default: edge_mask_reg_512p1[328] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101: edge_mask_reg_512p1[329] <= 1'b1;
 		default: edge_mask_reg_512p1[329] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101: edge_mask_reg_512p1[330] <= 1'b1;
 		default: edge_mask_reg_512p1[330] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000100,
12'b101000101,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001100010,
12'b11001100011: edge_mask_reg_512p1[331] <= 1'b1;
 		default: edge_mask_reg_512p1[331] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100: edge_mask_reg_512p1[332] <= 1'b1;
 		default: edge_mask_reg_512p1[332] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110000,
12'b10000110001,
12'b10000110011,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010010,
12'b11001010011,
12'b11001010100: edge_mask_reg_512p1[333] <= 1'b1;
 		default: edge_mask_reg_512p1[333] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110011,
12'b100110100,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110000,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110000,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10100110001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010010,
12'b11001010011,
12'b11001010100: edge_mask_reg_512p1[334] <= 1'b1;
 		default: edge_mask_reg_512p1[334] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110000,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b11001000011,
12'b11001000100: edge_mask_reg_512p1[335] <= 1'b1;
 		default: edge_mask_reg_512p1[335] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110011,
12'b110100,
12'b110101,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001011000,
12'b10001011001,
12'b10001101000,
12'b10001101001,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010011,
12'b10101010100,
12'b11001000011,
12'b11001000100: edge_mask_reg_512p1[336] <= 1'b1;
 		default: edge_mask_reg_512p1[336] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100100011,
12'b100100100,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b1000100011,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101101000,
12'b1101101001,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001011000,
12'b10001011001,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10101000011,
12'b10101000100: edge_mask_reg_512p1[337] <= 1'b1;
 		default: edge_mask_reg_512p1[337] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100100011,
12'b100100100,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101010100,
12'b1101010101,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101101000,
12'b1101101001,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10100110001,
12'b10100110011,
12'b10100110100,
12'b10101000011,
12'b10101000100: edge_mask_reg_512p1[338] <= 1'b1;
 		default: edge_mask_reg_512p1[338] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100011,
12'b100100,
12'b100101,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101011000,
12'b1101011001,
12'b10000100001,
12'b10000100010,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10100110011,
12'b10100110100: edge_mask_reg_512p1[339] <= 1'b1;
 		default: edge_mask_reg_512p1[339] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101011000,
12'b1101011001,
12'b10000100001,
12'b10000100010,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000011,
12'b10001000100: edge_mask_reg_512p1[340] <= 1'b1;
 		default: edge_mask_reg_512p1[340] <= 1'b0;
 	endcase

    case({x,y,z})
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101011000,
12'b1101011001,
12'b10000100100,
12'b10000110011,
12'b10000110100: edge_mask_reg_512p1[341] <= 1'b1;
 		default: edge_mask_reg_512p1[341] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001,
12'b10010,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100010001,
12'b100010010,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001001000,
12'b1001001001,
12'b1001011000,
12'b1001011001,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b10000100100,
12'b10000110011,
12'b10000110100: edge_mask_reg_512p1[342] <= 1'b1;
 		default: edge_mask_reg_512p1[342] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001,
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100010001,
12'b100010010,
12'b100010011,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001001000,
12'b1001001001,
12'b1001011000,
12'b1001011001,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100110011,
12'b1100110100,
12'b1100110101: edge_mask_reg_512p1[343] <= 1'b1;
 		default: edge_mask_reg_512p1[343] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b1000010010,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1100100100: edge_mask_reg_512p1[344] <= 1'b1;
 		default: edge_mask_reg_512p1[344] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101001000,
12'b101001001,
12'b101011000,
12'b101011001,
12'b1000100011,
12'b1000100100,
12'b1000100101: edge_mask_reg_512p1[345] <= 1'b1;
 		default: edge_mask_reg_512p1[345] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b100010010,
12'b100010100,
12'b100010101,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110100,
12'b100110101,
12'b101001000,
12'b101001001,
12'b101011000,
12'b101011001: edge_mask_reg_512p1[346] <= 1'b1;
 		default: edge_mask_reg_512p1[346] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110101,
12'b110110,
12'b110111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1011000,
12'b1011001,
12'b100010100,
12'b100010101,
12'b100100100,
12'b100100101: edge_mask_reg_512p1[347] <= 1'b1;
 		default: edge_mask_reg_512p1[347] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b10110,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b111010,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10011000,
12'b10011001,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100100111,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111000,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1000010010,
12'b1000010011,
12'b1000010100,
12'b1000010101,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000100110,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1000111000,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1100010010,
12'b1100010011,
12'b1100010100,
12'b1100010101,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100100110,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10000010010,
12'b10000010011,
12'b10000100010,
12'b10000100011,
12'b10000100100,
12'b10000100101,
12'b10000100110,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10000110111,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10100100010,
12'b10100100011,
12'b10100100100,
12'b10100100101,
12'b10100100110,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10100110110,
12'b10100110111,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101000111,
12'b10101001000,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101011010,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11000100010,
12'b11000100011,
12'b11000100100,
12'b11000100101,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11000110101,
12'b11000110110,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11100100010,
12'b11100100011,
12'b11100100100,
12'b11100100101,
12'b11100110010,
12'b11100110011,
12'b11100110100,
12'b11100110101,
12'b11100110110,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101000111,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100000100010,
12'b100000110010,
12'b100000110011,
12'b100000110100,
12'b100000110101,
12'b100000110110,
12'b100001000010,
12'b100001000011,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100100110010,
12'b100100110011,
12'b100100110100,
12'b100100110101,
12'b100101000010,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010010,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101000110010,
12'b101000110011,
12'b101001000010,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001010010,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101000010,
12'b101101000011,
12'b101101000100,
12'b101101000101,
12'b101101010010,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b110001010010,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110101010010,
12'b110101100010,
12'b110101100011,
12'b110101100100,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110110000010,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b111010000010: edge_mask_reg_512p1[348] <= 1'b1;
 		default: edge_mask_reg_512p1[348] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10011,
12'b10100,
12'b10101,
12'b100011,
12'b100100,
12'b100101,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1011000,
12'b1011001: edge_mask_reg_512p1[349] <= 1'b1;
 		default: edge_mask_reg_512p1[349] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100101100101,
12'b100101100110,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110110000010,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b111010000010: edge_mask_reg_512p1[350] <= 1'b1;
 		default: edge_mask_reg_512p1[350] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110101,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011: edge_mask_reg_512p1[351] <= 1'b1;
 		default: edge_mask_reg_512p1[351] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b100001100010,
12'b100001100011,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100101110001,
12'b100110000001: edge_mask_reg_512p1[352] <= 1'b1;
 		default: edge_mask_reg_512p1[352] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100101110001,
12'b100101110010,
12'b100110000001,
12'b100110000010: edge_mask_reg_512p1[353] <= 1'b1;
 		default: edge_mask_reg_512p1[353] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010010,
12'b100001010011,
12'b100001010100,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101100000,
12'b100101100001,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010100,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100010,
12'b110001100011,
12'b110001110010,
12'b110001110011: edge_mask_reg_512p1[354] <= 1'b1;
 		default: edge_mask_reg_512p1[354] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b11000110001,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11100110001,
12'b11100110010,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b100001000001,
12'b100001000010: edge_mask_reg_512p1[355] <= 1'b1;
 		default: edge_mask_reg_512p1[355] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110000,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101101000,
12'b10101101001,
12'b11000110001,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11100110001,
12'b11100110010,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b100001000001,
12'b100001000010: edge_mask_reg_512p1[356] <= 1'b1;
 		default: edge_mask_reg_512p1[356] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110011,
12'b100110100,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110000,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101101000,
12'b10101101001,
12'b11000110001,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11100110001,
12'b11100110010,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b100001000001,
12'b100001000010: edge_mask_reg_512p1[357] <= 1'b1;
 		default: edge_mask_reg_512p1[357] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001001,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101101000,
12'b10101101001,
12'b11000110001,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11100110001,
12'b11100110010,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b100001000001,
12'b100001000010: edge_mask_reg_512p1[358] <= 1'b1;
 		default: edge_mask_reg_512p1[358] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110011,
12'b110100,
12'b110101,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101001010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001000111,
12'b10001001001,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10100110001,
12'b10100110010,
12'b10100110011,
12'b10100110100,
12'b10100110101,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101000110,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101101000,
12'b10101101001,
12'b11000110001,
12'b11000110010,
12'b11000110011,
12'b11000110100,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001000101,
12'b11001000110,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11100110001,
12'b11100110010,
12'b11101000001,
12'b11101000010,
12'b11101000011,
12'b11101000100,
12'b11101000101,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b100001000001,
12'b100001000010: edge_mask_reg_512p1[359] <= 1'b1;
 		default: edge_mask_reg_512p1[359] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[360] <= 1'b1;
 		default: edge_mask_reg_512p1[360] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b10110110010,
12'b10110110011,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010110010,
12'b11010110011,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100: edge_mask_reg_512p1[361] <= 1'b1;
 		default: edge_mask_reg_512p1[361] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[362] <= 1'b1;
 		default: edge_mask_reg_512p1[362] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[363] <= 1'b1;
 		default: edge_mask_reg_512p1[363] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10,
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110101,
12'b110110,
12'b110111,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1011000,
12'b1011001,
12'b100010100,
12'b100010101,
12'b100100100,
12'b100100101: edge_mask_reg_512p1[364] <= 1'b1;
 		default: edge_mask_reg_512p1[364] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10,
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110101,
12'b110110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1011000,
12'b1011001,
12'b100010100,
12'b100010101,
12'b100100100,
12'b100100101: edge_mask_reg_512p1[365] <= 1'b1;
 		default: edge_mask_reg_512p1[365] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010110110,
12'b11010110111,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110011,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110100100,
12'b110110110100: edge_mask_reg_512p1[366] <= 1'b1;
 		default: edge_mask_reg_512p1[366] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010110110,
12'b11010110111,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110101,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110100,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110011,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p1[367] <= 1'b1;
 		default: edge_mask_reg_512p1[367] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100,
12'b10101,
12'b100100,
12'b100101,
12'b1001000,
12'b1001001,
12'b1011000,
12'b1011001: edge_mask_reg_512p1[368] <= 1'b1;
 		default: edge_mask_reg_512p1[368] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001,
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1001001000,
12'b1001001001,
12'b1001011000,
12'b1001011001,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100110011,
12'b1100110100,
12'b1100110101: edge_mask_reg_512p1[369] <= 1'b1;
 		default: edge_mask_reg_512p1[369] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001,
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b100010001,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b101000100,
12'b101000101,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1001001000: edge_mask_reg_512p1[370] <= 1'b1;
 		default: edge_mask_reg_512p1[370] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110110000101,
12'b110110000110,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110010110,
12'b110110100011,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b111010010011: edge_mask_reg_512p1[371] <= 1'b1;
 		default: edge_mask_reg_512p1[371] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110110,
12'b100110110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110110000101,
12'b110110000110,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110010110,
12'b110110100011,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101,
12'b111010010011: edge_mask_reg_512p1[372] <= 1'b1;
 		default: edge_mask_reg_512p1[372] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101100110,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b101001100110,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101001111000,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110010000010,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110101110110,
12'b110101110111,
12'b110110000010,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b110110000110,
12'b110110000111,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110010110,
12'b110110010111,
12'b111001110011,
12'b111001110100,
12'b111010000010,
12'b111010000011,
12'b111010000100,
12'b111010000101,
12'b111010010100,
12'b111010010101,
12'b111110000100: edge_mask_reg_512p1[373] <= 1'b1;
 		default: edge_mask_reg_512p1[373] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101110111,
12'b101111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[374] <= 1'b1;
 		default: edge_mask_reg_512p1[374] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101110111,
12'b101111000,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[375] <= 1'b1;
 		default: edge_mask_reg_512p1[375] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[376] <= 1'b1;
 		default: edge_mask_reg_512p1[376] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100010,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100101110010,
12'b100101110011,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100001,
12'b100110100010,
12'b101010000011,
12'b101010000100,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010100010: edge_mask_reg_512p1[377] <= 1'b1;
 		default: edge_mask_reg_512p1[377] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001011001,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101101001,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001000110,
12'b100001000111,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101000101,
12'b100101000110,
12'b100101000111,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101011000,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b101001000101,
12'b101001000110,
12'b101001000111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001011000,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101101000101,
12'b101101000110,
12'b101101000111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101100011,
12'b110101100100,
12'b110101100101,
12'b110101100110,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110101110110: edge_mask_reg_512p1[378] <= 1'b1;
 		default: edge_mask_reg_512p1[378] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111001001,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b1111010110,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000001,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011010001,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10011010101,
12'b10011010110,
12'b10011100011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111010010,
12'b10111010011,
12'b10111010100,
12'b10111010101,
12'b11011000101,
12'b11011010011: edge_mask_reg_512p1[379] <= 1'b1;
 		default: edge_mask_reg_512p1[379] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111001,
12'b1111000001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111010001,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b1111010110,
12'b1111100010,
12'b1111100011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10011010101,
12'b10011010110,
12'b10011100010,
12'b10011100011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111010010,
12'b10111010011,
12'b10111010100,
12'b10111010101,
12'b11011000101,
12'b11011010011: edge_mask_reg_512p1[380] <= 1'b1;
 		default: edge_mask_reg_512p1[380] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11001001,
12'b11001010,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11010101,
12'b11010110,
12'b11100001,
12'b11100010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111100001,
12'b111100010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000001,
12'b1011000010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011010001,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1011100010,
12'b1011100011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111001,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b1111010110,
12'b1111100010,
12'b1111100011,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10011010101,
12'b10011010110,
12'b10011100010,
12'b10011100011,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111010010,
12'b10111010011,
12'b10111010100,
12'b10111010101,
12'b11011000101,
12'b11011010011: edge_mask_reg_512p1[381] <= 1'b1;
 		default: edge_mask_reg_512p1[381] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100001,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100010010,
12'b100010011,
12'b100100001,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111000,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b1000100001,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1100100001,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100110001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101011000,
12'b1101011001,
12'b10000100001,
12'b10000100010,
12'b10000100011,
12'b10000100100,
12'b10000100101,
12'b10000110001,
12'b10000110010,
12'b10000110011,
12'b10000110100,
12'b10000110101,
12'b10000110110,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10100110011,
12'b10100110100,
12'b10100110101: edge_mask_reg_512p1[382] <= 1'b1;
 		default: edge_mask_reg_512p1[382] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1101110010,
12'b1101110011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001101000,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110011000,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010010000,
12'b100010010001: edge_mask_reg_512p1[383] <= 1'b1;
 		default: edge_mask_reg_512p1[383] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10100110,
12'b10100111,
12'b10101000,
12'b10110100,
12'b10110101,
12'b10110110,
12'b10110111,
12'b10111000,
12'b11000000,
12'b11000001,
12'b11000010,
12'b11000011,
12'b11000100,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11010000,
12'b11010001,
12'b11010010,
12'b11010011,
12'b11010100,
12'b11100010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110110110,
12'b110110111,
12'b110111000,
12'b111000001,
12'b111000010,
12'b111000011,
12'b111000100,
12'b111000101,
12'b111010000,
12'b111010001,
12'b111010010,
12'b111010011,
12'b111010100,
12'b1011010010,
12'b1011010011: edge_mask_reg_512p1[384] <= 1'b1;
 		default: edge_mask_reg_512p1[384] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110010,
12'b1110011,
12'b1110100,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100010,
12'b101100011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110000,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110100,
12'b101110101,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010010,
12'b110010011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010101,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[385] <= 1'b1;
 		default: edge_mask_reg_512p1[385] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010000,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101110010001,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100001,
12'b101110100010: edge_mask_reg_512p1[386] <= 1'b1;
 		default: edge_mask_reg_512p1[386] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000000,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010010,
12'b10010011,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[387] <= 1'b1;
 		default: edge_mask_reg_512p1[387] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[388] <= 1'b1;
 		default: edge_mask_reg_512p1[388] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[389] <= 1'b1;
 		default: edge_mask_reg_512p1[389] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b100001110111,
12'b100001111000,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100101110110,
12'b100101110111,
12'b100101111000,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110001000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100110,
12'b100110100111,
12'b101001110110,
12'b101001110111,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010001000,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101101110110,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110000111,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b110001110110,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010000111,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b110110000110,
12'b110110000111,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110010110,
12'b110110010111,
12'b111010010011,
12'b111010010100: edge_mask_reg_512p1[390] <= 1'b1;
 		default: edge_mask_reg_512p1[390] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110010010,
12'b11110010011,
12'b11110010100: edge_mask_reg_512p1[391] <= 1'b1;
 		default: edge_mask_reg_512p1[391] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100000,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110101000,
12'b10110101001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000011,
12'b11110000100,
12'b11110010010,
12'b11110010011,
12'b11110010100: edge_mask_reg_512p1[392] <= 1'b1;
 		default: edge_mask_reg_512p1[392] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[393] <= 1'b1;
 		default: edge_mask_reg_512p1[393] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[394] <= 1'b1;
 		default: edge_mask_reg_512p1[394] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110011,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001100010,
12'b11001100011: edge_mask_reg_512p1[395] <= 1'b1;
 		default: edge_mask_reg_512p1[395] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110011,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100: edge_mask_reg_512p1[396] <= 1'b1;
 		default: edge_mask_reg_512p1[396] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000111,
12'b10110001000,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010111,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[397] <= 1'b1;
 		default: edge_mask_reg_512p1[397] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000111,
12'b10110001000,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010111,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010010,
12'b11101010011,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[398] <= 1'b1;
 		default: edge_mask_reg_512p1[398] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110010,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100001,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110110010: edge_mask_reg_512p1[399] <= 1'b1;
 		default: edge_mask_reg_512p1[399] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110010,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100001,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110110010: edge_mask_reg_512p1[400] <= 1'b1;
 		default: edge_mask_reg_512p1[400] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110010,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010110010,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100001,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110110010,
12'b110010100010: edge_mask_reg_512p1[401] <= 1'b1;
 		default: edge_mask_reg_512p1[401] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010100001,
12'b100010100011,
12'b100010100100,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[402] <= 1'b1;
 		default: edge_mask_reg_512p1[402] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110100010,
12'b11110100011,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100: edge_mask_reg_512p1[403] <= 1'b1;
 		default: edge_mask_reg_512p1[403] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110110000,
12'b11110110001,
12'b11110110010,
12'b11110110011: edge_mask_reg_512p1[404] <= 1'b1;
 		default: edge_mask_reg_512p1[404] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b10110110110,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11010110100,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110110000,
12'b11110110001,
12'b11110110010,
12'b11110110011: edge_mask_reg_512p1[405] <= 1'b1;
 		default: edge_mask_reg_512p1[405] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010000,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100000,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[406] <= 1'b1;
 		default: edge_mask_reg_512p1[406] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010000,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100000,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10110111,
12'b10111000,
12'b10111001,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100001,
12'b110100010,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[407] <= 1'b1;
 		default: edge_mask_reg_512p1[407] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[408] <= 1'b1;
 		default: edge_mask_reg_512p1[408] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[409] <= 1'b1;
 		default: edge_mask_reg_512p1[409] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110111000,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[410] <= 1'b1;
 		default: edge_mask_reg_512p1[410] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101011000,
12'b1101011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010010,
12'b100110010011,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101110000001,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b101110010010,
12'b101110010011,
12'b110010000010,
12'b110010000011: edge_mask_reg_512p1[411] <= 1'b1;
 		default: edge_mask_reg_512p1[411] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110010,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110010,
12'b101010110011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110100001,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110110010,
12'b101110110011,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100010,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011,
12'b110110010011,
12'b110110010100,
12'b110110100011,
12'b110110100100: edge_mask_reg_512p1[412] <= 1'b1;
 		default: edge_mask_reg_512p1[412] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110010,
12'b1110110011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110010,
12'b10110110011,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[413] <= 1'b1;
 		default: edge_mask_reg_512p1[413] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010101000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[414] <= 1'b1;
 		default: edge_mask_reg_512p1[414] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110000,
12'b11010110001,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[415] <= 1'b1;
 		default: edge_mask_reg_512p1[415] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110110,
12'b101001110101,
12'b101001110110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101101110100,
12'b101101110101,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010010,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011,
12'b110010110100,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b110110010010,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110100011,
12'b110110100100: edge_mask_reg_512p1[416] <= 1'b1;
 		default: edge_mask_reg_512p1[416] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b100001110110,
12'b100001110111,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010001000,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100101110110,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110000111,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b101001110101,
12'b101001110110,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010000111,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010110011,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101101110100,
12'b101101110101,
12'b101110000011,
12'b101110000100,
12'b101110000101,
12'b101110000110,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110011,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b110010000011,
12'b110010000100,
12'b110010000101,
12'b110010000110,
12'b110010010010,
12'b110010010011,
12'b110010010100,
12'b110010010101,
12'b110010010110,
12'b110010100011,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010110011,
12'b110010110100,
12'b110110000011,
12'b110110000100,
12'b110110000101,
12'b110110010010,
12'b110110010011,
12'b110110010100,
12'b110110010101,
12'b110110100011,
12'b110110100100,
12'b110110110100: edge_mask_reg_512p1[417] <= 1'b1;
 		default: edge_mask_reg_512p1[417] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101110000100,
12'b101110000101,
12'b101110010001,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b110010010010: edge_mask_reg_512p1[418] <= 1'b1;
 		default: edge_mask_reg_512p1[418] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001111000,
12'b11001111001,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010000110,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101110000100,
12'b101110000101,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b110010010010: edge_mask_reg_512p1[419] <= 1'b1;
 		default: edge_mask_reg_512p1[419] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11110000111,
12'b11110001000,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[420] <= 1'b1;
 		default: edge_mask_reg_512p1[420] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10010,
12'b10011,
12'b10100,
12'b10101,
12'b100010,
12'b100011,
12'b100100,
12'b100101,
12'b100110,
12'b100111,
12'b110011,
12'b110100,
12'b110101,
12'b110110,
12'b110111,
12'b111000,
12'b111001,
12'b111010,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1001011,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b100010010,
12'b100010011,
12'b100010100,
12'b100010101,
12'b100100010,
12'b100100011,
12'b100100100,
12'b100100101,
12'b100100110,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100110101,
12'b100110110,
12'b100110111,
12'b100111000,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101101001,
12'b1000010010,
12'b1000010011,
12'b1000100010,
12'b1000100011,
12'b1000100100,
12'b1000100101,
12'b1000100110,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1000110101,
12'b1000110110,
12'b1000110111,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1100100010,
12'b1100100011,
12'b1100100100,
12'b1100100101,
12'b1100100110,
12'b1100110011,
12'b1100110100,
12'b1100110101,
12'b1100110110,
12'b1100110111,
12'b10000100100,
12'b10000100101,
12'b10000110100,
12'b10000110101: edge_mask_reg_512p1[421] <= 1'b1;
 		default: edge_mask_reg_512p1[421] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[422] <= 1'b1;
 		default: edge_mask_reg_512p1[422] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110101000,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[423] <= 1'b1;
 		default: edge_mask_reg_512p1[423] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000000,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010010,
12'b10010011,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100111,
12'b1010101000,
12'b1101110010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11110000111,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[424] <= 1'b1;
 		default: edge_mask_reg_512p1[424] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001000111,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101000110,
12'b10101000111,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110011,
12'b101101110100,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[425] <= 1'b1;
 		default: edge_mask_reg_512p1[425] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110011,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010000,
12'b100110010001,
12'b100110010010,
12'b100110010011: edge_mask_reg_512p1[426] <= 1'b1;
 		default: edge_mask_reg_512p1[426] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010101000,
12'b1010101001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b1110101001,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10010101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11101110011,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100010,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010100001,
12'b100010100010,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010000,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110100001,
12'b100110100010,
12'b101010000011,
12'b101010000100,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010100010: edge_mask_reg_512p1[427] <= 1'b1;
 		default: edge_mask_reg_512p1[427] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010: edge_mask_reg_512p1[428] <= 1'b1;
 		default: edge_mask_reg_512p1[428] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000100,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000001,
12'b100110000010,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010,
12'b101101110001,
12'b101101110010: edge_mask_reg_512p1[429] <= 1'b1;
 		default: edge_mask_reg_512p1[429] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001101000,
12'b11001101001,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010011000,
12'b11010011001,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010001,
12'b100110010010,
12'b101001110011,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010010001: edge_mask_reg_512p1[430] <= 1'b1;
 		default: edge_mask_reg_512p1[430] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010110111,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000100,
12'b101111000101,
12'b110010010101,
12'b110010010110,
12'b110010010111,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110011000100,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p1[431] <= 1'b1;
 		default: edge_mask_reg_512p1[431] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111001,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100111,
12'b11010101000,
12'b11010101001,
12'b11010110111,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110011001,
12'b11110100110,
12'b11110100111,
12'b11110101000,
12'b11110101001,
12'b11110110110,
12'b11110110111,
12'b11110111000,
12'b100010010110,
12'b100010010111,
12'b100010011000,
12'b100010100110,
12'b100010100111,
12'b100010101000,
12'b100010110110,
12'b100010110111,
12'b100010111000,
12'b100110010110,
12'b100110010111,
12'b100110011000,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110101000,
12'b100110110101,
12'b100110110110,
12'b100110110111,
12'b100110111000,
12'b101010010101,
12'b101010010110,
12'b101010010111,
12'b101010011000,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010100111,
12'b101010101000,
12'b101010110100,
12'b101010110101,
12'b101010110110,
12'b101010110111,
12'b101010111000,
12'b101110010101,
12'b101110010110,
12'b101110010111,
12'b101110100100,
12'b101110100101,
12'b101110100110,
12'b101110100111,
12'b101110110100,
12'b101110110101,
12'b101110110110,
12'b101110110111,
12'b101111000100,
12'b101111000101,
12'b110010010110,
12'b110010010111,
12'b110010100100,
12'b110010100101,
12'b110010100110,
12'b110010100111,
12'b110010110100,
12'b110010110101,
12'b110010110110,
12'b110010110111,
12'b110011000100,
12'b110110100100,
12'b110110100101,
12'b110110110100,
12'b110110110101: edge_mask_reg_512p1[432] <= 1'b1;
 		default: edge_mask_reg_512p1[432] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010100,
12'b101010101,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100101,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110001000,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010001000,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011,
12'b11101110010,
12'b11101110011: edge_mask_reg_512p1[433] <= 1'b1;
 		default: edge_mask_reg_512p1[433] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010100,
12'b101010101,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100101,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101100010,
12'b11101100011: edge_mask_reg_512p1[434] <= 1'b1;
 		default: edge_mask_reg_512p1[434] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010100,
12'b101010101,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100101,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100000,
12'b1001100001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001010010,
12'b11001010011,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010001000,
12'b11101100010,
12'b11101100011,
12'b11101110010,
12'b11101110011,
12'b11101110100: edge_mask_reg_512p1[435] <= 1'b1;
 		default: edge_mask_reg_512p1[435] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110010000,
12'b100110010001,
12'b100110010010: edge_mask_reg_512p1[436] <= 1'b1;
 		default: edge_mask_reg_512p1[436] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110100111,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110010110,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[437] <= 1'b1;
 		default: edge_mask_reg_512p1[437] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010001,
12'b100010000001: edge_mask_reg_512p1[438] <= 1'b1;
 		default: edge_mask_reg_512p1[438] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100010,
12'b1101100011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010001,
12'b100010000001: edge_mask_reg_512p1[439] <= 1'b1;
 		default: edge_mask_reg_512p1[439] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000100,
12'b1010000101,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001101000,
12'b10001101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b101010000001,
12'b101010000010,
12'b101010010001,
12'b101010010010: edge_mask_reg_512p1[440] <= 1'b1;
 		default: edge_mask_reg_512p1[440] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010011000,
12'b11010011001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b101010000001,
12'b101010000010,
12'b101010010001,
12'b101010010010: edge_mask_reg_512p1[441] <= 1'b1;
 		default: edge_mask_reg_512p1[441] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110101010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011001,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010010011,
12'b100010010100: edge_mask_reg_512p1[442] <= 1'b1;
 		default: edge_mask_reg_512p1[442] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10101011,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b10111010,
12'b11000101,
12'b11000110,
12'b11000111,
12'b11001000,
12'b11010101,
12'b11010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b110111010,
12'b111000100,
12'b111000101,
12'b111000110,
12'b111000111,
12'b111001000,
12'b111010100,
12'b111010101,
12'b111010110,
12'b111010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1010111010,
12'b1011000011,
12'b1011000100,
12'b1011000101,
12'b1011000110,
12'b1011000111,
12'b1011001000,
12'b1011010010,
12'b1011010011,
12'b1011010100,
12'b1011010101,
12'b1011010110,
12'b1011010111,
12'b1011100101,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1111000010,
12'b1111000011,
12'b1111000100,
12'b1111000101,
12'b1111000110,
12'b1111000111,
12'b1111010010,
12'b1111010011,
12'b1111010100,
12'b1111010101,
12'b1111010110,
12'b1111100010,
12'b1111100011,
12'b1111100100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10011000010,
12'b10011000011,
12'b10011000100,
12'b10011000101,
12'b10011000110,
12'b10011000111,
12'b10011010010,
12'b10011010011,
12'b10011010100,
12'b10011010101,
12'b10011010110,
12'b10011100011,
12'b10011100100,
12'b10111000011,
12'b10111000100,
12'b10111000101,
12'b10111000110,
12'b10111010010,
12'b10111010011,
12'b10111010100,
12'b10111010101,
12'b10111010110,
12'b10111100011,
12'b10111100100,
12'b11011000101,
12'b11011010011,
12'b11011010100,
12'b11011100011: edge_mask_reg_512p1[443] <= 1'b1;
 		default: edge_mask_reg_512p1[443] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[444] <= 1'b1;
 		default: edge_mask_reg_512p1[444] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[445] <= 1'b1;
 		default: edge_mask_reg_512p1[445] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[446] <= 1'b1;
 		default: edge_mask_reg_512p1[446] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100010,
12'b1001100011,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110000,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[447] <= 1'b1;
 		default: edge_mask_reg_512p1[447] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010001011,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010011000,
12'b11010011001,
12'b11101110000,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110001000,
12'b11110001001,
12'b11110010001,
12'b100010000001: edge_mask_reg_512p1[448] <= 1'b1;
 		default: edge_mask_reg_512p1[448] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10001011,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10011011,
12'b10101000,
12'b10101001,
12'b10101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110101000,
12'b110101001,
12'b110101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010011011,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11010101000,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110011000,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b11110110011,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100010100111,
12'b100010110010,
12'b100010110011,
12'b100010110100,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110100111,
12'b100110110010,
12'b100110110011,
12'b100110110100,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110011,
12'b101010110100,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110110011: edge_mask_reg_512p1[449] <= 1'b1;
 		default: edge_mask_reg_512p1[449] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000000,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[450] <= 1'b1;
 		default: edge_mask_reg_512p1[450] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000000,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[451] <= 1'b1;
 		default: edge_mask_reg_512p1[451] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000000,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[452] <= 1'b1;
 		default: edge_mask_reg_512p1[452] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001111000,
12'b11001111001,
12'b11101000000,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100010,
12'b11101100011,
12'b11101100100: edge_mask_reg_512p1[453] <= 1'b1;
 		default: edge_mask_reg_512p1[453] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101111000,
12'b10101111001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100011: edge_mask_reg_512p1[454] <= 1'b1;
 		default: edge_mask_reg_512p1[454] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11101000001,
12'b11101000010,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100: edge_mask_reg_512p1[455] <= 1'b1;
 		default: edge_mask_reg_512p1[455] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000100,
12'b101000101,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11101000001,
12'b11101000010,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100: edge_mask_reg_512p1[456] <= 1'b1;
 		default: edge_mask_reg_512p1[456] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110010,
12'b1000110011,
12'b1000110100,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1100110010,
12'b1100110011,
12'b1100110100,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b10000110000,
12'b10000110001,
12'b10000110011,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001000110,
12'b10001001000,
12'b10001001001,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001111000,
12'b10001111001,
12'b10101000000,
12'b10101000001,
12'b10101000010,
12'b10101000011,
12'b10101000100,
12'b10101000101,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101101000,
12'b10101101001,
12'b11001000000,
12'b11001000001,
12'b11001000010,
12'b11001000011,
12'b11001000100,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11101000001,
12'b11101000010,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100: edge_mask_reg_512p1[457] <= 1'b1;
 		default: edge_mask_reg_512p1[457] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b10110110101,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110010,
12'b11010110011,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[458] <= 1'b1;
 		default: edge_mask_reg_512p1[458] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010111000,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110010,
12'b11010110011: edge_mask_reg_512p1[459] <= 1'b1;
 		default: edge_mask_reg_512p1[459] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110001011,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010011010,
12'b11010100101,
12'b11010100110,
12'b11010100111,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b11110100111,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110010111,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b100110100110,
12'b100110110010,
12'b100110110011,
12'b101010000100,
12'b101010000101,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101010100110,
12'b101010110010,
12'b101010110011,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b101110100100,
12'b101110100101,
12'b101110110010,
12'b101110110011,
12'b110010100010,
12'b110010100011: edge_mask_reg_512p1[460] <= 1'b1;
 		default: edge_mask_reg_512p1[460] <= 1'b0;
 	endcase

    case({x,y,z})
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100110,
12'b10100111,
12'b10101000,
12'b10101001,
12'b10101010,
12'b10110110,
12'b10110111,
12'b10111000,
12'b10111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100000,
12'b110100011,
12'b110100100,
12'b110100101,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110000,
12'b110110011,
12'b110110100,
12'b110110101,
12'b110110110,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100000,
12'b1010100001,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110000,
12'b1010110001,
12'b1010110010,
12'b1010110011,
12'b1010110100,
12'b1010110101,
12'b1010110110,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110000,
12'b1110110001,
12'b1110110010,
12'b1110110011,
12'b1110110100,
12'b1110110101,
12'b1110110110,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10010000111,
12'b10010001000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010110000,
12'b10010110001,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10010110101,
12'b10010110110,
12'b10010110111,
12'b10010111000,
12'b10010111001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100111,
12'b10110101000,
12'b10110110000,
12'b10110110001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010010010,
12'b11010010011,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010110010,
12'b11010110011: edge_mask_reg_512p1[461] <= 1'b1;
 		default: edge_mask_reg_512p1[461] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000000,
12'b10000001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000101,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010000,
12'b10010001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010101,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10100110,
12'b10100111,
12'b10101000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110001,
12'b1101110010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110010100,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010101000,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[462] <= 1'b1;
 		default: edge_mask_reg_512p1[462] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110010,
12'b1001110011,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110011000: edge_mask_reg_512p1[463] <= 1'b1;
 		default: edge_mask_reg_512p1[463] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110011000: edge_mask_reg_512p1[464] <= 1'b1;
 		default: edge_mask_reg_512p1[464] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[465] <= 1'b1;
 		default: edge_mask_reg_512p1[465] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110011,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010111,
12'b11010011000,
12'b11110000111,
12'b11110001000,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[466] <= 1'b1;
 		default: edge_mask_reg_512p1[466] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000000,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[467] <= 1'b1;
 		default: edge_mask_reg_512p1[467] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000010,
12'b10000011,
12'b10000100,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010010,
12'b10010011,
12'b10010100,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000111,
12'b11110001000,
12'b11110011000: edge_mask_reg_512p1[468] <= 1'b1;
 		default: edge_mask_reg_512p1[468] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[469] <= 1'b1;
 		default: edge_mask_reg_512p1[469] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100010,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10101010010,
12'b10101010011,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101101000,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100: edge_mask_reg_512p1[470] <= 1'b1;
 		default: edge_mask_reg_512p1[470] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011001,
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100011,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100000,
12'b1101100001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101101000,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000010,
12'b11110000011,
12'b11110000100: edge_mask_reg_512p1[471] <= 1'b1;
 		default: edge_mask_reg_512p1[471] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[472] <= 1'b1;
 		default: edge_mask_reg_512p1[472] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[473] <= 1'b1;
 		default: edge_mask_reg_512p1[473] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[474] <= 1'b1;
 		default: edge_mask_reg_512p1[474] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110001000,
12'b11110001001: edge_mask_reg_512p1[475] <= 1'b1;
 		default: edge_mask_reg_512p1[475] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011: edge_mask_reg_512p1[476] <= 1'b1;
 		default: edge_mask_reg_512p1[476] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100: edge_mask_reg_512p1[477] <= 1'b1;
 		default: edge_mask_reg_512p1[477] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100110,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100: edge_mask_reg_512p1[478] <= 1'b1;
 		default: edge_mask_reg_512p1[478] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100100,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101001000,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110010,
12'b11001110011,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b100001010000,
12'b100001010001,
12'b100001010011,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011: edge_mask_reg_512p1[479] <= 1'b1;
 		default: edge_mask_reg_512p1[479] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1010111,
12'b1011000,
12'b1011001,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100101,
12'b1001100110,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1101001000,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b10001010000,
12'b10001010001,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100000,
12'b10001100001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10101000010,
12'b10101000011,
12'b10101010000,
12'b10101010001,
12'b10101010010,
12'b10101010011,
12'b10101010100,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100000,
12'b10101100001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b11001000010,
12'b11001000011,
12'b11001010000,
12'b11001010001,
12'b11001010010,
12'b11001010011,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001011000,
12'b11001100000,
12'b11001100001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010000,
12'b11101010001,
12'b11101010010,
12'b11101010011,
12'b11101010100,
12'b11101100000,
12'b11101100001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b100001010000,
12'b100001010001,
12'b100001010011,
12'b100001100000,
12'b100001100001,
12'b100001100010,
12'b100001100011: edge_mask_reg_512p1[480] <= 1'b1;
 		default: edge_mask_reg_512p1[480] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110110111,
12'b110111000,
12'b110111001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010110111,
12'b1010111000,
12'b1010111001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110001011,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110011011,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b1110110011,
12'b1110110111,
12'b1110111000,
12'b1110111001,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10010110010,
12'b10010110011,
12'b10010110100,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110100111,
12'b10110101000,
12'b10110101001,
12'b10110110010,
12'b10110110011,
12'b10110110100,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11010101000,
12'b11010110010,
12'b11010110011,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100110010001: edge_mask_reg_512p1[481] <= 1'b1;
 		default: edge_mask_reg_512p1[481] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1101000,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001101000,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[482] <= 1'b1;
 		default: edge_mask_reg_512p1[482] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101101000,
12'b1101101001,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[483] <= 1'b1;
 		default: edge_mask_reg_512p1[483] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100110,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110010,
12'b101110011,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000010,
12'b110000011,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000000,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[484] <= 1'b1;
 		default: edge_mask_reg_512p1[484] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010110,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110110,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110010,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101110000,
12'b1101110001,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110101000,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001110000,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010101000,
12'b10101100100,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[485] <= 1'b1;
 		default: edge_mask_reg_512p1[485] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110011,
12'b101001110100,
12'b101001110110,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110011,
12'b101101110100,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[486] <= 1'b1;
 		default: edge_mask_reg_512p1[486] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110110,
12'b100101110111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110011,
12'b101001110100,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110011,
12'b101101110100,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001110011,
12'b110101100011,
12'b110101100100: edge_mask_reg_512p1[487] <= 1'b1;
 		default: edge_mask_reg_512p1[487] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1011011,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101011011,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001011011,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101011011,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001000111,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101000110,
12'b10101000111,
12'b10101010101,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001001,
12'b10110001010,
12'b11001000101,
12'b11001000110,
12'b11001000111,
12'b11001010100,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11101000100,
12'b11101000101,
12'b11101000110,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b100001000100,
12'b100001000101,
12'b100001000110,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101000011,
12'b100101000100,
12'b100101000101,
12'b100101000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b101001000011,
12'b101001000100,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001110011,
12'b101001110100,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110011,
12'b110001010011,
12'b110001010100,
12'b110001100011,
12'b110001100100: edge_mask_reg_512p1[488] <= 1'b1;
 		default: edge_mask_reg_512p1[488] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[489] <= 1'b1;
 		default: edge_mask_reg_512p1[489] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[490] <= 1'b1;
 		default: edge_mask_reg_512p1[490] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[491] <= 1'b1;
 		default: edge_mask_reg_512p1[491] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[492] <= 1'b1;
 		default: edge_mask_reg_512p1[492] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110000,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000000,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[493] <= 1'b1;
 		default: edge_mask_reg_512p1[493] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[494] <= 1'b1;
 		default: edge_mask_reg_512p1[494] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100: edge_mask_reg_512p1[495] <= 1'b1;
 		default: edge_mask_reg_512p1[495] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001000,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100101100011,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b101001110001,
12'b101010000001: edge_mask_reg_512p1[496] <= 1'b1;
 		default: edge_mask_reg_512p1[496] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b10001100101,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010001010,
12'b11010011000,
12'b11010011001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b11101111001,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110001001,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100010000000,
12'b100010000001,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101100011,
12'b100101100100,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100: edge_mask_reg_512p1[497] <= 1'b1;
 		default: edge_mask_reg_512p1[497] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10001010,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10011010,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110011011,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010011011,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10010101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11001111000,
12'b11001111001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010110,
12'b11010010111,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010100110,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b11110010000,
12'b11110010001,
12'b11110010010,
12'b11110010011,
12'b11110010100,
12'b11110010101,
12'b11110010110,
12'b11110010111,
12'b11110100000,
12'b11110100001,
12'b11110100010,
12'b11110100011,
12'b11110100100,
12'b11110100101,
12'b11110100110,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100010000111,
12'b100010010000,
12'b100010010001,
12'b100010010010,
12'b100010010011,
12'b100010010100,
12'b100010010101,
12'b100010010110,
12'b100010010111,
12'b100010100000,
12'b100010100001,
12'b100010100010,
12'b100010100011,
12'b100010100100,
12'b100010100101,
12'b100010100110,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110010001,
12'b100110010010,
12'b100110010011,
12'b100110010100,
12'b100110010101,
12'b100110010110,
12'b100110100001,
12'b100110100010,
12'b100110100011,
12'b100110100100,
12'b100110100101,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101010010001,
12'b101010010010,
12'b101010010011,
12'b101010010100,
12'b101010010101,
12'b101010010110,
12'b101010100001,
12'b101010100010,
12'b101010100011,
12'b101010100100,
12'b101010100101,
12'b101110010010,
12'b101110010011,
12'b101110010100,
12'b101110010101,
12'b101110100010,
12'b101110100011,
12'b101110100100: edge_mask_reg_512p1[498] <= 1'b1;
 		default: edge_mask_reg_512p1[498] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010001011,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001010101,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11110000101,
12'b11110000110,
12'b11110000111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110010,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100010000010,
12'b100010000011,
12'b100010000100,
12'b100010000101,
12'b100010000110,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110001,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100110000001,
12'b100110000010,
12'b100110000011,
12'b100110000100,
12'b100110000101,
12'b100110000110,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101010000001,
12'b101010000010,
12'b101010000011,
12'b101010000100,
12'b101010000101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101110000010,
12'b101110000011,
12'b101110000100,
12'b110001100010,
12'b110001100011,
12'b110001110010,
12'b110001110011,
12'b110010000010: edge_mask_reg_512p1[499] <= 1'b1;
 		default: edge_mask_reg_512p1[499] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[500] <= 1'b1;
 		default: edge_mask_reg_512p1[500] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b10010111,
12'b10011000,
12'b10011001,
12'b10100111,
12'b10101000,
12'b10101001,
12'b101110111,
12'b101111000,
12'b101111001,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110010100,
12'b110010101,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110011010,
12'b110100111,
12'b110101000,
12'b110101001,
12'b110101010,
12'b110111000,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100010,
12'b1010100011,
12'b1010100100,
12'b1010100101,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1010101010,
12'b1010111000,
12'b1010111001,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100001,
12'b1110100010,
12'b1110100011,
12'b1110100100,
12'b1110100101,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b1110101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100001,
12'b10010100010,
12'b10010100011,
12'b10010100100,
12'b10010100101,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100001,
12'b10110100010,
12'b10110100011,
12'b10110100100,
12'b10110100101,
12'b10110100110,
12'b10110101000,
12'b10110101001,
12'b11010000010,
12'b11010000011,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010011000,
12'b11010011001,
12'b11010100000,
12'b11010100001,
12'b11010100010,
12'b11010100011,
12'b11010100100,
12'b11010100101,
12'b11010101000,
12'b11110010010,
12'b11110010011,
12'b11110100010,
12'b11110100011: edge_mask_reg_512p1[501] <= 1'b1;
 		default: edge_mask_reg_512p1[501] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110111,
12'b1111000,
12'b1111001,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110011,
12'b1001110100,
12'b1001110101,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000011,
12'b1010000100,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101100011,
12'b1101100100,
12'b1101100101,
12'b1101100110,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110010,
12'b1101110011,
12'b1101110100,
12'b1101110101,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110011000,
12'b1110011001,
12'b10001100010,
12'b10001100011,
12'b10001100100,
12'b10001100101,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010011000,
12'b10010011001,
12'b10101100010,
12'b10101100011,
12'b10101100100,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110000,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110011000,
12'b10110011001,
12'b11001100010,
12'b11001100011,
12'b11001100100,
12'b11001100101,
12'b11001101000,
12'b11001101001,
12'b11001110000,
12'b11001110001,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010001000,
12'b11010001001,
12'b11101100010,
12'b11101100011,
12'b11101100100,
12'b11101110000,
12'b11101110001,
12'b11101110010,
12'b11101110011,
12'b11101110100,
12'b11101110101,
12'b11101111000,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b100001110000,
12'b100001110001,
12'b100001110010,
12'b100010000000,
12'b100010000001: edge_mask_reg_512p1[502] <= 1'b1;
 		default: edge_mask_reg_512p1[502] <= 1'b0;
 	endcase

    case({x,y,z})
12'b110000,
12'b110001,
12'b110010,
12'b110011,
12'b110100,
12'b110101,
12'b111000,
12'b111001,
12'b1000000,
12'b1000001,
12'b1000010,
12'b1000011,
12'b1000100,
12'b1000101,
12'b1000110,
12'b1000111,
12'b1001000,
12'b1001001,
12'b1001010,
12'b1010010,
12'b1010011,
12'b1010100,
12'b1010101,
12'b1010110,
12'b1010111,
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b100110000,
12'b100110001,
12'b100110010,
12'b100110011,
12'b100110100,
12'b100111000,
12'b101000000,
12'b101000001,
12'b101000010,
12'b101000011,
12'b101000100,
12'b101000101,
12'b101000110,
12'b101000111,
12'b101001000,
12'b101001001,
12'b101001010,
12'b101010000,
12'b101010001,
12'b101010010,
12'b101010011,
12'b101010100,
12'b101010101,
12'b101010110,
12'b101010111,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b1000110000,
12'b1000110001,
12'b1000110010,
12'b1000110011,
12'b1001000000,
12'b1001000001,
12'b1001000010,
12'b1001000011,
12'b1001000100,
12'b1001000101,
12'b1001000110,
12'b1001000111,
12'b1001001000,
12'b1001001001,
12'b1001010000,
12'b1001010001,
12'b1001010010,
12'b1001010011,
12'b1001010100,
12'b1001010101,
12'b1001010110,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1101000000,
12'b1101000001,
12'b1101000010,
12'b1101000011,
12'b1101000100,
12'b1101000101,
12'b1101000110,
12'b1101000111,
12'b1101001000,
12'b1101001001,
12'b1101010000,
12'b1101010001,
12'b1101010010,
12'b1101010011,
12'b1101010100,
12'b1101010101,
12'b1101010110,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b10001000000,
12'b10001000001,
12'b10001000010,
12'b10001000011,
12'b10001000100,
12'b10001000101,
12'b10001010010,
12'b10001010011,
12'b10001010100,
12'b10001010101,
12'b10001010110,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10101000011,
12'b10101010010,
12'b10101010011: edge_mask_reg_512p1[503] <= 1'b1;
 		default: edge_mask_reg_512p1[503] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b1111011,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101101011,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1101111011,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101011001,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010001001,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101011000,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110111,
12'b11101111000,
12'b100001000110,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001011000,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100001111000,
12'b100101000101,
12'b100101000110,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b101001000101,
12'b101001000110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001010111,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110110,
12'b101001110111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101010111,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001010111,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110001110111,
12'b110101010011,
12'b110101010100,
12'b110101010101,
12'b110101010110,
12'b110101100011,
12'b110101100100,
12'b110101100101,
12'b110101100110,
12'b110101100111,
12'b110101110011,
12'b110101110100,
12'b110101110110,
12'b111001010011,
12'b111001010100,
12'b111001100011,
12'b111001100100,
12'b111001100101: edge_mask_reg_512p1[504] <= 1'b1;
 		default: edge_mask_reg_512p1[504] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010100,
12'b101001010101,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010100,
12'b101101010101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110101100010,
12'b110101100011,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b111001110010,
12'b111001110011: edge_mask_reg_512p1[505] <= 1'b1;
 		default: edge_mask_reg_512p1[505] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010100,
12'b101101010101,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110101100010,
12'b110101100011,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b111001110010,
12'b111001110011: edge_mask_reg_512p1[506] <= 1'b1;
 		default: edge_mask_reg_512p1[506] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1011000,
12'b1011001,
12'b1011010,
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1101011,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b110001010,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001101011,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10001111011,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101010110,
12'b10101010111,
12'b10101011000,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001010111,
12'b11001011000,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010101,
12'b11101010110,
12'b11101010111,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010100,
12'b100001010101,
12'b100001010110,
12'b100001010111,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001101000,
12'b100001110110,
12'b100001110111,
12'b100101010100,
12'b100101010101,
12'b100101010110,
12'b100101010111,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101101000,
12'b100101110110,
12'b100101110111,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001010110,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001100111,
12'b101001101000,
12'b101001110101,
12'b101001110110,
12'b101001110111,
12'b101101010011,
12'b101101010100,
12'b101101010101,
12'b101101010110,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101100111,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b101101110111,
12'b110001010011,
12'b110001010100,
12'b110001010101,
12'b110001010110,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001100110,
12'b110001100111,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110001110110,
12'b110101010011,
12'b110101010100,
12'b110101100011,
12'b110101100100,
12'b110101100101,
12'b110101100110,
12'b110101100111,
12'b110101110011,
12'b110101110100,
12'b110101110101,
12'b110101110110,
12'b111001100011,
12'b111001100100,
12'b111001100101,
12'b111001110100: edge_mask_reg_512p1[507] <= 1'b1;
 		default: edge_mask_reg_512p1[507] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100001,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001110010,
12'b110001110011: edge_mask_reg_512p1[508] <= 1'b1;
 		default: edge_mask_reg_512p1[508] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1101010,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101011001,
12'b101011010,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101101011,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b101111011,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001011010,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001101011,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1001111011,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101011010,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001011010,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b11001010101,
12'b11001010110,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001101010,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11001111010,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101010110,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101101000,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b100001010011,
12'b100001010100,
12'b100001010101,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101010101,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b101001010011,
12'b101001010100,
12'b101001010101,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101010100,
12'b101101010101,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b110001100001,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110101100010,
12'b110101100011: edge_mask_reg_512p1[509] <= 1'b1;
 		default: edge_mask_reg_512p1[509] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1100111,
12'b1101000,
12'b1101001,
12'b1110110,
12'b1110111,
12'b1111000,
12'b1111001,
12'b1111010,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10001001,
12'b101011000,
12'b101100111,
12'b101101000,
12'b101101001,
12'b101101010,
12'b101110111,
12'b101111000,
12'b101111001,
12'b101111010,
12'b110000111,
12'b110001000,
12'b110001001,
12'b1001010111,
12'b1001011000,
12'b1001011001,
12'b1001100111,
12'b1001101000,
12'b1001101001,
12'b1001101010,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1001111010,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1101010111,
12'b1101011000,
12'b1101011001,
12'b1101100111,
12'b1101101000,
12'b1101101001,
12'b1101101010,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b10001010111,
12'b10001011000,
12'b10001011001,
12'b10001100110,
12'b10001100111,
12'b10001101000,
12'b10001101001,
12'b10001101010,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10101011000,
12'b10101011001,
12'b10101100101,
12'b10101100110,
12'b10101100111,
12'b10101101000,
12'b10101101001,
12'b10101101010,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10101111010,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b11001100100,
12'b11001100101,
12'b11001100110,
12'b11001100111,
12'b11001101000,
12'b11001101001,
12'b11001110100,
12'b11001110101,
12'b11001110110,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010001000,
12'b11010001001,
12'b11101010011,
12'b11101010100,
12'b11101010101,
12'b11101100011,
12'b11101100100,
12'b11101100101,
12'b11101100110,
12'b11101100111,
12'b11101110100,
12'b11101110101,
12'b11101110110,
12'b11101110111,
12'b11101111000,
12'b100001010011,
12'b100001010100,
12'b100001100010,
12'b100001100011,
12'b100001100100,
12'b100001100101,
12'b100001100110,
12'b100001100111,
12'b100001110011,
12'b100001110100,
12'b100001110101,
12'b100001110110,
12'b100001110111,
12'b100101010011,
12'b100101010100,
12'b100101100010,
12'b100101100011,
12'b100101100100,
12'b100101100101,
12'b100101100110,
12'b100101100111,
12'b100101110010,
12'b100101110011,
12'b100101110100,
12'b100101110101,
12'b100101110110,
12'b100101110111,
12'b101001010011,
12'b101001010100,
12'b101001100001,
12'b101001100010,
12'b101001100011,
12'b101001100100,
12'b101001100101,
12'b101001100110,
12'b101001110001,
12'b101001110010,
12'b101001110011,
12'b101001110100,
12'b101001110101,
12'b101001110110,
12'b101101100001,
12'b101101100010,
12'b101101100011,
12'b101101100100,
12'b101101100101,
12'b101101100110,
12'b101101110001,
12'b101101110010,
12'b101101110011,
12'b101101110100,
12'b101101110101,
12'b101101110110,
12'b110001100001,
12'b110001100010,
12'b110001100011,
12'b110001100100,
12'b110001100101,
12'b110001110010,
12'b110001110011,
12'b110001110100,
12'b110001110101,
12'b110010000010,
12'b110010000011,
12'b110101100010,
12'b110101100011,
12'b110101110010,
12'b110101110011,
12'b110101110100,
12'b111001110010,
12'b111001110011: edge_mask_reg_512p1[510] <= 1'b1;
 		default: edge_mask_reg_512p1[510] <= 1'b0;
 	endcase

    case({x,y,z})
12'b1110110,
12'b1110111,
12'b1111000,
12'b10000110,
12'b10000111,
12'b10001000,
12'b10010110,
12'b10010111,
12'b10011000,
12'b101110110,
12'b101110111,
12'b101111000,
12'b110000001,
12'b110000010,
12'b110000011,
12'b110000100,
12'b110000101,
12'b110000110,
12'b110000111,
12'b110001000,
12'b110010001,
12'b110010010,
12'b110010011,
12'b110010100,
12'b110010110,
12'b110010111,
12'b110011000,
12'b110011001,
12'b110100110,
12'b110100111,
12'b110101000,
12'b110101001,
12'b1001110110,
12'b1001110111,
12'b1001111000,
12'b1001111001,
12'b1010000001,
12'b1010000010,
12'b1010000011,
12'b1010000100,
12'b1010000101,
12'b1010000110,
12'b1010000111,
12'b1010001000,
12'b1010001001,
12'b1010001010,
12'b1010010000,
12'b1010010001,
12'b1010010010,
12'b1010010011,
12'b1010010100,
12'b1010010101,
12'b1010010110,
12'b1010010111,
12'b1010011000,
12'b1010011001,
12'b1010011010,
12'b1010100110,
12'b1010100111,
12'b1010101000,
12'b1010101001,
12'b1101110110,
12'b1101110111,
12'b1101111000,
12'b1101111001,
12'b1101111010,
12'b1110000000,
12'b1110000001,
12'b1110000010,
12'b1110000011,
12'b1110000100,
12'b1110000101,
12'b1110000110,
12'b1110000111,
12'b1110001000,
12'b1110001001,
12'b1110001010,
12'b1110010000,
12'b1110010001,
12'b1110010010,
12'b1110010011,
12'b1110010100,
12'b1110010101,
12'b1110010110,
12'b1110010111,
12'b1110011000,
12'b1110011001,
12'b1110011010,
12'b1110100000,
12'b1110100110,
12'b1110100111,
12'b1110101000,
12'b1110101001,
12'b10001110010,
12'b10001110011,
12'b10001110100,
12'b10001110101,
12'b10001110110,
12'b10001110111,
12'b10001111000,
12'b10001111001,
12'b10001111010,
12'b10010000000,
12'b10010000001,
12'b10010000010,
12'b10010000011,
12'b10010000100,
12'b10010000101,
12'b10010000110,
12'b10010000111,
12'b10010001000,
12'b10010001001,
12'b10010001010,
12'b10010010000,
12'b10010010001,
12'b10010010010,
12'b10010010011,
12'b10010010100,
12'b10010010101,
12'b10010010110,
12'b10010010111,
12'b10010011000,
12'b10010011001,
12'b10010011010,
12'b10010100000,
12'b10010100110,
12'b10010100111,
12'b10010101000,
12'b10010101001,
12'b10101110001,
12'b10101110010,
12'b10101110011,
12'b10101110100,
12'b10101110101,
12'b10101110110,
12'b10101110111,
12'b10101111000,
12'b10101111001,
12'b10110000000,
12'b10110000001,
12'b10110000010,
12'b10110000011,
12'b10110000100,
12'b10110000101,
12'b10110000110,
12'b10110000111,
12'b10110001000,
12'b10110001001,
12'b10110001010,
12'b10110010000,
12'b10110010001,
12'b10110010010,
12'b10110010011,
12'b10110010100,
12'b10110010101,
12'b10110010110,
12'b10110010111,
12'b10110011000,
12'b10110011001,
12'b10110011010,
12'b10110100000,
12'b10110100111,
12'b10110101000,
12'b11001110010,
12'b11001110011,
12'b11001110100,
12'b11001110111,
12'b11001111000,
12'b11001111001,
12'b11010000000,
12'b11010000001,
12'b11010000010,
12'b11010000011,
12'b11010000100,
12'b11010000101,
12'b11010000110,
12'b11010000111,
12'b11010001000,
12'b11010001001,
12'b11010010000,
12'b11010010001,
12'b11010010010,
12'b11010010011,
12'b11010010100,
12'b11010010101,
12'b11010010111,
12'b11010011000,
12'b11101110010,
12'b11101110011,
12'b11110000000,
12'b11110000001,
12'b11110000010,
12'b11110000011,
12'b11110000100,
12'b11110000111,
12'b11110001000,
12'b11110010000,
12'b11110010001,
12'b11110010111,
12'b11110011000: edge_mask_reg_512p1[511] <= 1'b1;
 		default: edge_mask_reg_512p1[511] <= 1'b0;
 	endcase

end
endmodule

