/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 7
second: 18
********************************************/

module prm_LUTX1_Ca_3_4_4_chk512p4(
	input [2:0] x,
	input [3:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p4
);

	reg [511:0] edge_mask_reg_512p4;
	assign edge_mask_512p4= edge_mask_reg_512p4;

always @( *) begin
    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101100011,
11'b1101100100,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[0] <= 1'b1;
 		default: edge_mask_reg_512p4[0] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101000111,
11'b101001000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1101010111,
11'b1101011000,
11'b1101100111,
11'b1101101000,
11'b1101110111,
11'b1101111000: edge_mask_reg_512p4[1] <= 1'b1;
 		default: edge_mask_reg_512p4[1] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[2] <= 1'b1;
 		default: edge_mask_reg_512p4[2] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100110,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p4[3] <= 1'b1;
 		default: edge_mask_reg_512p4[3] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11101110100,
11'b11101110101,
11'b11110000011,
11'b11110000100,
11'b11110000101,
11'b11110010011,
11'b11110010100: edge_mask_reg_512p4[4] <= 1'b1;
 		default: edge_mask_reg_512p4[4] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11100010,
11'b111010001,
11'b111010010,
11'b111010011: edge_mask_reg_512p4[5] <= 1'b1;
 		default: edge_mask_reg_512p4[5] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110111000,
11'b110111001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100001,
11'b10010100010: edge_mask_reg_512p4[6] <= 1'b1;
 		default: edge_mask_reg_512p4[6] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10010000000,
11'b10010000001,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p4[7] <= 1'b1;
 		default: edge_mask_reg_512p4[7] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10110110100,
11'b10110110101,
11'b10110110110: edge_mask_reg_512p4[8] <= 1'b1;
 		default: edge_mask_reg_512p4[8] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100110,
11'b1101100111,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001100101,
11'b11001100110,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100,
11'b11110000101,
11'b11110010011,
11'b11110010100: edge_mask_reg_512p4[9] <= 1'b1;
 		default: edge_mask_reg_512p4[9] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p4[10] <= 1'b1;
 		default: edge_mask_reg_512p4[10] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110110000,
11'b1110110001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[11] <= 1'b1;
 		default: edge_mask_reg_512p4[11] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b1001000011,
11'b1001000100,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1101000011,
11'b1101000100,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100: edge_mask_reg_512p4[12] <= 1'b1;
 		default: edge_mask_reg_512p4[12] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[13] <= 1'b1;
 		default: edge_mask_reg_512p4[13] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11001000,
11'b11010011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110100011,
11'b1110100100,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[14] <= 1'b1;
 		default: edge_mask_reg_512p4[14] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110000,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000000,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[15] <= 1'b1;
 		default: edge_mask_reg_512p4[15] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000011,
11'b10011000100,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b11010010110,
11'b11010010111,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110011,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000100,
11'b11011000101,
11'b11110110101: edge_mask_reg_512p4[16] <= 1'b1;
 		default: edge_mask_reg_512p4[16] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p4[17] <= 1'b1;
 		default: edge_mask_reg_512p4[17] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[18] <= 1'b1;
 		default: edge_mask_reg_512p4[18] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[19] <= 1'b1;
 		default: edge_mask_reg_512p4[19] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110010,
11'b10001110011,
11'b10010000010,
11'b10010000011,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[20] <= 1'b1;
 		default: edge_mask_reg_512p4[20] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100011,
11'b10010100100,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101: edge_mask_reg_512p4[21] <= 1'b1;
 		default: edge_mask_reg_512p4[21] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[22] <= 1'b1;
 		default: edge_mask_reg_512p4[22] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[23] <= 1'b1;
 		default: edge_mask_reg_512p4[23] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100: edge_mask_reg_512p4[24] <= 1'b1;
 		default: edge_mask_reg_512p4[24] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b11001000011,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11101000100,
11'b11101000101,
11'b11101010100,
11'b11101010101: edge_mask_reg_512p4[25] <= 1'b1;
 		default: edge_mask_reg_512p4[25] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[26] <= 1'b1;
 		default: edge_mask_reg_512p4[26] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[27] <= 1'b1;
 		default: edge_mask_reg_512p4[27] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[28] <= 1'b1;
 		default: edge_mask_reg_512p4[28] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[29] <= 1'b1;
 		default: edge_mask_reg_512p4[29] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[30] <= 1'b1;
 		default: edge_mask_reg_512p4[30] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[31] <= 1'b1;
 		default: edge_mask_reg_512p4[31] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[32] <= 1'b1;
 		default: edge_mask_reg_512p4[32] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[33] <= 1'b1;
 		default: edge_mask_reg_512p4[33] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[34] <= 1'b1;
 		default: edge_mask_reg_512p4[34] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[35] <= 1'b1;
 		default: edge_mask_reg_512p4[35] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[36] <= 1'b1;
 		default: edge_mask_reg_512p4[36] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[37] <= 1'b1;
 		default: edge_mask_reg_512p4[37] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[38] <= 1'b1;
 		default: edge_mask_reg_512p4[38] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[39] <= 1'b1;
 		default: edge_mask_reg_512p4[39] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[40] <= 1'b1;
 		default: edge_mask_reg_512p4[40] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[41] <= 1'b1;
 		default: edge_mask_reg_512p4[41] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[42] <= 1'b1;
 		default: edge_mask_reg_512p4[42] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[43] <= 1'b1;
 		default: edge_mask_reg_512p4[43] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[44] <= 1'b1;
 		default: edge_mask_reg_512p4[44] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[45] <= 1'b1;
 		default: edge_mask_reg_512p4[45] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[46] <= 1'b1;
 		default: edge_mask_reg_512p4[46] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[47] <= 1'b1;
 		default: edge_mask_reg_512p4[47] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b10101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[48] <= 1'b1;
 		default: edge_mask_reg_512p4[48] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[49] <= 1'b1;
 		default: edge_mask_reg_512p4[49] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[50] <= 1'b1;
 		default: edge_mask_reg_512p4[50] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[51] <= 1'b1;
 		default: edge_mask_reg_512p4[51] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101100101,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b10001100011,
11'b10001100100,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[52] <= 1'b1;
 		default: edge_mask_reg_512p4[52] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100101,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10001100011,
11'b10001100100,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11010000010,
11'b11010000011,
11'b11010010011: edge_mask_reg_512p4[53] <= 1'b1;
 		default: edge_mask_reg_512p4[53] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11110011,
11'b11110100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111110011,
11'b111110100,
11'b1011010101,
11'b1011010110: edge_mask_reg_512p4[54] <= 1'b1;
 		default: edge_mask_reg_512p4[54] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11110011,
11'b11110100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111100111,
11'b111110011,
11'b111110100,
11'b1011000101,
11'b1011000110,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011100011,
11'b1011100100,
11'b1011100101,
11'b1011100110: edge_mask_reg_512p4[55] <= 1'b1;
 		default: edge_mask_reg_512p4[55] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[56] <= 1'b1;
 		default: edge_mask_reg_512p4[56] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p4[57] <= 1'b1;
 		default: edge_mask_reg_512p4[57] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10001110001,
11'b10001110010,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000: edge_mask_reg_512p4[58] <= 1'b1;
 		default: edge_mask_reg_512p4[58] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110001000,
11'b1110001001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10101100001,
11'b10101100010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[59] <= 1'b1;
 		default: edge_mask_reg_512p4[59] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[60] <= 1'b1;
 		default: edge_mask_reg_512p4[60] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101: edge_mask_reg_512p4[61] <= 1'b1;
 		default: edge_mask_reg_512p4[61] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110010001,
11'b10110010010,
11'b10110100010: edge_mask_reg_512p4[62] <= 1'b1;
 		default: edge_mask_reg_512p4[62] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[63] <= 1'b1;
 		default: edge_mask_reg_512p4[63] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010: edge_mask_reg_512p4[64] <= 1'b1;
 		default: edge_mask_reg_512p4[64] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[65] <= 1'b1;
 		default: edge_mask_reg_512p4[65] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[66] <= 1'b1;
 		default: edge_mask_reg_512p4[66] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b10001110011,
11'b10001110100,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010: edge_mask_reg_512p4[67] <= 1'b1;
 		default: edge_mask_reg_512p4[67] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100: edge_mask_reg_512p4[68] <= 1'b1;
 		default: edge_mask_reg_512p4[68] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101: edge_mask_reg_512p4[69] <= 1'b1;
 		default: edge_mask_reg_512p4[69] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010100,
11'b11101110100,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[70] <= 1'b1;
 		default: edge_mask_reg_512p4[70] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100011,
11'b11001100100,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010100,
11'b11101110100,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[71] <= 1'b1;
 		default: edge_mask_reg_512p4[71] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b111010101,
11'b111010110: edge_mask_reg_512p4[72] <= 1'b1;
 		default: edge_mask_reg_512p4[72] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010111,
11'b101011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1101100001,
11'b1101100010,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[73] <= 1'b1;
 		default: edge_mask_reg_512p4[73] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[74] <= 1'b1;
 		default: edge_mask_reg_512p4[74] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[75] <= 1'b1;
 		default: edge_mask_reg_512p4[75] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[76] <= 1'b1;
 		default: edge_mask_reg_512p4[76] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b101101000,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[77] <= 1'b1;
 		default: edge_mask_reg_512p4[77] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[78] <= 1'b1;
 		default: edge_mask_reg_512p4[78] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10101000,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[79] <= 1'b1;
 		default: edge_mask_reg_512p4[79] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110110111,
11'b110111000,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111010010,
11'b111010011: edge_mask_reg_512p4[80] <= 1'b1;
 		default: edge_mask_reg_512p4[80] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[81] <= 1'b1;
 		default: edge_mask_reg_512p4[81] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10101000010,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b11001000100,
11'b11001000101,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111: edge_mask_reg_512p4[82] <= 1'b1;
 		default: edge_mask_reg_512p4[82] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110010,
11'b10001110011,
11'b10101010000,
11'b10101010001,
11'b10101100000,
11'b10101100001: edge_mask_reg_512p4[83] <= 1'b1;
 		default: edge_mask_reg_512p4[83] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11,
11'b100,
11'b101,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110101,
11'b110110,
11'b110111,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100010100,
11'b100010101: edge_mask_reg_512p4[84] <= 1'b1;
 		default: edge_mask_reg_512p4[84] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000010,
11'b10010010100,
11'b10010010101,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[85] <= 1'b1;
 		default: edge_mask_reg_512p4[85] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000010,
11'b1011000011,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000010,
11'b1111000011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10110110011,
11'b10110110100: edge_mask_reg_512p4[86] <= 1'b1;
 		default: edge_mask_reg_512p4[86] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10110100011,
11'b10110110011: edge_mask_reg_512p4[87] <= 1'b1;
 		default: edge_mask_reg_512p4[87] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001010100,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010100,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001001,
11'b1110001010,
11'b10001100010,
11'b10001100011,
11'b10001110010,
11'b10001110011,
11'b10010000010: edge_mask_reg_512p4[88] <= 1'b1;
 		default: edge_mask_reg_512p4[88] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[89] <= 1'b1;
 		default: edge_mask_reg_512p4[89] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10110100011,
11'b10110100100: edge_mask_reg_512p4[90] <= 1'b1;
 		default: edge_mask_reg_512p4[90] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010101001,
11'b1010101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10001110100,
11'b10001110101,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[91] <= 1'b1;
 		default: edge_mask_reg_512p4[91] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10110010011,
11'b10110010100,
11'b10110100011: edge_mask_reg_512p4[92] <= 1'b1;
 		default: edge_mask_reg_512p4[92] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b1111100,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[93] <= 1'b1;
 		default: edge_mask_reg_512p4[93] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[94] <= 1'b1;
 		default: edge_mask_reg_512p4[94] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[95] <= 1'b1;
 		default: edge_mask_reg_512p4[95] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[96] <= 1'b1;
 		default: edge_mask_reg_512p4[96] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[97] <= 1'b1;
 		default: edge_mask_reg_512p4[97] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[98] <= 1'b1;
 		default: edge_mask_reg_512p4[98] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100010,
11'b11100011,
11'b11100100,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[99] <= 1'b1;
 		default: edge_mask_reg_512p4[99] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[100] <= 1'b1;
 		default: edge_mask_reg_512p4[100] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[101] <= 1'b1;
 		default: edge_mask_reg_512p4[101] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101001000,
11'b101001001,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101111000,
11'b1101111001,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10101000010,
11'b10101000011,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101100001,
11'b10101100010: edge_mask_reg_512p4[102] <= 1'b1;
 		default: edge_mask_reg_512p4[102] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10110010110,
11'b10110010111,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000100,
11'b11011000101,
11'b11011000110: edge_mask_reg_512p4[103] <= 1'b1;
 		default: edge_mask_reg_512p4[103] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[104] <= 1'b1;
 		default: edge_mask_reg_512p4[104] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b11001000100,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100100,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p4[105] <= 1'b1;
 		default: edge_mask_reg_512p4[105] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001011001,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100100,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p4[106] <= 1'b1;
 		default: edge_mask_reg_512p4[106] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11,
11'b100,
11'b101,
11'b110,
11'b111,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b10111,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1101001,
11'b100000011,
11'b100000100,
11'b100000101,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100010111,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111: edge_mask_reg_512p4[107] <= 1'b1;
 		default: edge_mask_reg_512p4[107] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1101110010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[108] <= 1'b1;
 		default: edge_mask_reg_512p4[108] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[109] <= 1'b1;
 		default: edge_mask_reg_512p4[109] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010: edge_mask_reg_512p4[110] <= 1'b1;
 		default: edge_mask_reg_512p4[110] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011: edge_mask_reg_512p4[111] <= 1'b1;
 		default: edge_mask_reg_512p4[111] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010011,
11'b110010100,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1011000001,
11'b1011000010: edge_mask_reg_512p4[112] <= 1'b1;
 		default: edge_mask_reg_512p4[112] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010100100: edge_mask_reg_512p4[113] <= 1'b1;
 		default: edge_mask_reg_512p4[113] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000001: edge_mask_reg_512p4[114] <= 1'b1;
 		default: edge_mask_reg_512p4[114] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110011,
11'b1110110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110100000,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[115] <= 1'b1;
 		default: edge_mask_reg_512p4[115] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001111000,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110011,
11'b1110110100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110100000,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[116] <= 1'b1;
 		default: edge_mask_reg_512p4[116] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110: edge_mask_reg_512p4[117] <= 1'b1;
 		default: edge_mask_reg_512p4[117] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100010,
11'b10010100011: edge_mask_reg_512p4[118] <= 1'b1;
 		default: edge_mask_reg_512p4[118] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110001,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11101010010,
11'b11101010011,
11'b11101100010,
11'b11101100011,
11'b11101110010,
11'b11101110011: edge_mask_reg_512p4[119] <= 1'b1;
 		default: edge_mask_reg_512p4[119] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110001,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11101110010,
11'b11101110011: edge_mask_reg_512p4[120] <= 1'b1;
 		default: edge_mask_reg_512p4[120] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000010,
11'b10011000011: edge_mask_reg_512p4[121] <= 1'b1;
 		default: edge_mask_reg_512p4[121] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10011000011,
11'b10011000100: edge_mask_reg_512p4[122] <= 1'b1;
 		default: edge_mask_reg_512p4[122] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011010011,
11'b1011010100,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111010011,
11'b10010100100,
11'b10010110100,
11'b10011000011: edge_mask_reg_512p4[123] <= 1'b1;
 		default: edge_mask_reg_512p4[123] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11110011,
11'b11110100,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100010,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111110011,
11'b111110100,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011100010,
11'b1011100011,
11'b1011100100,
11'b1011100101: edge_mask_reg_512p4[124] <= 1'b1;
 		default: edge_mask_reg_512p4[124] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010: edge_mask_reg_512p4[125] <= 1'b1;
 		default: edge_mask_reg_512p4[125] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110: edge_mask_reg_512p4[126] <= 1'b1;
 		default: edge_mask_reg_512p4[126] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100110011,
11'b100110100,
11'b100110101,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b10001000001,
11'b10001000010: edge_mask_reg_512p4[127] <= 1'b1;
 		default: edge_mask_reg_512p4[127] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000110011,
11'b1000110100,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010011,
11'b10001010100: edge_mask_reg_512p4[128] <= 1'b1;
 		default: edge_mask_reg_512p4[128] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011000,
11'b10011001,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010010,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010010,
11'b11001110010,
11'b11001110011,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p4[129] <= 1'b1;
 		default: edge_mask_reg_512p4[129] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b111000110,
11'b111000111,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111100110: edge_mask_reg_512p4[130] <= 1'b1;
 		default: edge_mask_reg_512p4[130] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[131] <= 1'b1;
 		default: edge_mask_reg_512p4[131] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[132] <= 1'b1;
 		default: edge_mask_reg_512p4[132] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[133] <= 1'b1;
 		default: edge_mask_reg_512p4[133] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000010,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[134] <= 1'b1;
 		default: edge_mask_reg_512p4[134] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b10010000010,
11'b10010000011,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[135] <= 1'b1;
 		default: edge_mask_reg_512p4[135] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b10010000010,
11'b10010000011,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[136] <= 1'b1;
 		default: edge_mask_reg_512p4[136] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b10010000010,
11'b10010000011,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[137] <= 1'b1;
 		default: edge_mask_reg_512p4[137] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010101001,
11'b1010101010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11010010011,
11'b11010010100,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p4[138] <= 1'b1;
 		default: edge_mask_reg_512p4[138] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101: edge_mask_reg_512p4[139] <= 1'b1;
 		default: edge_mask_reg_512p4[139] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[140] <= 1'b1;
 		default: edge_mask_reg_512p4[140] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110110,
11'b110111,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100010011,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b10000100010,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110010,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100100011,
11'b10100100100,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110: edge_mask_reg_512p4[141] <= 1'b1;
 		default: edge_mask_reg_512p4[141] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11110001,
11'b11110010,
11'b11110011,
11'b11110100,
11'b110100111,
11'b110101000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111100001,
11'b111100010,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111110001,
11'b111110010,
11'b111110011,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1011100001,
11'b1011100010,
11'b1011100011,
11'b1011100100,
11'b1011100101: edge_mask_reg_512p4[142] <= 1'b1;
 		default: edge_mask_reg_512p4[142] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b11100011,
11'b11100100,
11'b110111000,
11'b111000001,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111100011,
11'b111100100: edge_mask_reg_512p4[143] <= 1'b1;
 		default: edge_mask_reg_512p4[143] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11101110011,
11'b11101110100,
11'b11110000011,
11'b11110000100: edge_mask_reg_512p4[144] <= 1'b1;
 		default: edge_mask_reg_512p4[144] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101: edge_mask_reg_512p4[145] <= 1'b1;
 		default: edge_mask_reg_512p4[145] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101: edge_mask_reg_512p4[146] <= 1'b1;
 		default: edge_mask_reg_512p4[146] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101: edge_mask_reg_512p4[147] <= 1'b1;
 		default: edge_mask_reg_512p4[147] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101011000,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001: edge_mask_reg_512p4[148] <= 1'b1;
 		default: edge_mask_reg_512p4[148] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000: edge_mask_reg_512p4[149] <= 1'b1;
 		default: edge_mask_reg_512p4[149] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b11001110010,
11'b11001110011,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010011,
11'b11010010100: edge_mask_reg_512p4[150] <= 1'b1;
 		default: edge_mask_reg_512p4[150] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101: edge_mask_reg_512p4[151] <= 1'b1;
 		default: edge_mask_reg_512p4[151] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10101110011,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110011,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011: edge_mask_reg_512p4[152] <= 1'b1;
 		default: edge_mask_reg_512p4[152] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10101110011,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110011,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p4[153] <= 1'b1;
 		default: edge_mask_reg_512p4[153] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110011,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010001,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011: edge_mask_reg_512p4[154] <= 1'b1;
 		default: edge_mask_reg_512p4[154] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010110,
11'b11001010111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000011,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[155] <= 1'b1;
 		default: edge_mask_reg_512p4[155] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110001000,
11'b1110001001,
11'b10001110001,
11'b10001110010,
11'b10010000001: edge_mask_reg_512p4[156] <= 1'b1;
 		default: edge_mask_reg_512p4[156] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[157] <= 1'b1;
 		default: edge_mask_reg_512p4[157] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[158] <= 1'b1;
 		default: edge_mask_reg_512p4[158] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010: edge_mask_reg_512p4[159] <= 1'b1;
 		default: edge_mask_reg_512p4[159] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[160] <= 1'b1;
 		default: edge_mask_reg_512p4[160] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010011,
11'b11010100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111010001,
11'b1111010010,
11'b1111010011,
11'b1111010100: edge_mask_reg_512p4[161] <= 1'b1;
 		default: edge_mask_reg_512p4[161] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100000,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b110000,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1101000,
11'b1101001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100110010,
11'b100110011,
11'b100110100,
11'b101001000,
11'b101001001,
11'b101011000,
11'b101011001: edge_mask_reg_512p4[162] <= 1'b1;
 		default: edge_mask_reg_512p4[162] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10110000100,
11'b10110000101,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110011: edge_mask_reg_512p4[163] <= 1'b1;
 		default: edge_mask_reg_512p4[163] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110: edge_mask_reg_512p4[164] <= 1'b1;
 		default: edge_mask_reg_512p4[164] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011: edge_mask_reg_512p4[165] <= 1'b1;
 		default: edge_mask_reg_512p4[165] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[166] <= 1'b1;
 		default: edge_mask_reg_512p4[166] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011010011,
11'b1011010100: edge_mask_reg_512p4[167] <= 1'b1;
 		default: edge_mask_reg_512p4[167] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b11100011,
11'b11100100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011010011,
11'b1011010100: edge_mask_reg_512p4[168] <= 1'b1;
 		default: edge_mask_reg_512p4[168] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101: edge_mask_reg_512p4[169] <= 1'b1;
 		default: edge_mask_reg_512p4[169] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110101,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1011000,
11'b1011001: edge_mask_reg_512p4[170] <= 1'b1;
 		default: edge_mask_reg_512p4[170] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p4[171] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110010001,
11'b10110010010,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[172] <= 1'b1;
 		default: edge_mask_reg_512p4[172] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110010001,
11'b10110010010,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[173] <= 1'b1;
 		default: edge_mask_reg_512p4[173] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100001,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b10000110011,
11'b10000110101,
11'b10001000101: edge_mask_reg_512p4[174] <= 1'b1;
 		default: edge_mask_reg_512p4[174] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[175] <= 1'b1;
 		default: edge_mask_reg_512p4[175] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001110000,
11'b10001110001,
11'b10001110010: edge_mask_reg_512p4[176] <= 1'b1;
 		default: edge_mask_reg_512p4[176] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110001,
11'b10001110010: edge_mask_reg_512p4[177] <= 1'b1;
 		default: edge_mask_reg_512p4[177] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110000,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101101000: edge_mask_reg_512p4[178] <= 1'b1;
 		default: edge_mask_reg_512p4[178] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101010011,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110001,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100: edge_mask_reg_512p4[179] <= 1'b1;
 		default: edge_mask_reg_512p4[179] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010100,
11'b1101010101,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010100,
11'b10001010101,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[180] <= 1'b1;
 		default: edge_mask_reg_512p4[180] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11110100,
11'b11110101,
11'b11110110,
11'b11110111,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111100111,
11'b111110100,
11'b111110101,
11'b111110110: edge_mask_reg_512p4[181] <= 1'b1;
 		default: edge_mask_reg_512p4[181] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11110011,
11'b11110100,
11'b11110101,
11'b11110110,
11'b11110111: edge_mask_reg_512p4[182] <= 1'b1;
 		default: edge_mask_reg_512p4[182] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111010101,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10110110100,
11'b10110110101: edge_mask_reg_512p4[183] <= 1'b1;
 		default: edge_mask_reg_512p4[183] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100011: edge_mask_reg_512p4[184] <= 1'b1;
 		default: edge_mask_reg_512p4[184] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10001110011,
11'b10001110100,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[185] <= 1'b1;
 		default: edge_mask_reg_512p4[185] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p4[186] <= 1'b1;
 		default: edge_mask_reg_512p4[186] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10,
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100010100,
11'b100010101,
11'b100100011,
11'b100100100,
11'b100100101: edge_mask_reg_512p4[187] <= 1'b1;
 		default: edge_mask_reg_512p4[187] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10,
11'b11,
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100010010,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110: edge_mask_reg_512p4[188] <= 1'b1;
 		default: edge_mask_reg_512p4[188] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110101,
11'b100110110: edge_mask_reg_512p4[189] <= 1'b1;
 		default: edge_mask_reg_512p4[189] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[190] <= 1'b1;
 		default: edge_mask_reg_512p4[190] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[191] <= 1'b1;
 		default: edge_mask_reg_512p4[191] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11,
11'b100,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100000011,
11'b100000100,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001001,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[192] <= 1'b1;
 		default: edge_mask_reg_512p4[192] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100010,
11'b1101100011: edge_mask_reg_512p4[193] <= 1'b1;
 		default: edge_mask_reg_512p4[193] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[194] <= 1'b1;
 		default: edge_mask_reg_512p4[194] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101010011,
11'b10101010100,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001110001,
11'b11001110010: edge_mask_reg_512p4[195] <= 1'b1;
 		default: edge_mask_reg_512p4[195] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101110000,
11'b10101110001,
11'b10101110011,
11'b10110000000,
11'b10110000001,
11'b10110000011: edge_mask_reg_512p4[196] <= 1'b1;
 		default: edge_mask_reg_512p4[196] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010010111,
11'b1010011000,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1110110010,
11'b1110110011: edge_mask_reg_512p4[197] <= 1'b1;
 		default: edge_mask_reg_512p4[197] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10110000010: edge_mask_reg_512p4[198] <= 1'b1;
 		default: edge_mask_reg_512p4[198] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110111,
11'b1010111000: edge_mask_reg_512p4[199] <= 1'b1;
 		default: edge_mask_reg_512p4[199] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b11001110010: edge_mask_reg_512p4[200] <= 1'b1;
 		default: edge_mask_reg_512p4[200] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101110001,
11'b10101110011,
11'b10110000001: edge_mask_reg_512p4[201] <= 1'b1;
 		default: edge_mask_reg_512p4[201] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100011,
11'b100100,
11'b100101,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001011000,
11'b1001011001,
11'b1001101000,
11'b1001101001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1101000011,
11'b1101000100: edge_mask_reg_512p4[202] <= 1'b1;
 		default: edge_mask_reg_512p4[202] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[203] <= 1'b1;
 		default: edge_mask_reg_512p4[203] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10110110010,
11'b10110110011: edge_mask_reg_512p4[204] <= 1'b1;
 		default: edge_mask_reg_512p4[204] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110111,
11'b10111000,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p4[205] <= 1'b1;
 		default: edge_mask_reg_512p4[205] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101: edge_mask_reg_512p4[206] <= 1'b1;
 		default: edge_mask_reg_512p4[206] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101: edge_mask_reg_512p4[207] <= 1'b1;
 		default: edge_mask_reg_512p4[207] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000: edge_mask_reg_512p4[208] <= 1'b1;
 		default: edge_mask_reg_512p4[208] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010010,
11'b10110010011,
11'b11001110010,
11'b11001110011,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p4[209] <= 1'b1;
 		default: edge_mask_reg_512p4[209] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110011,
11'b110111000,
11'b110111001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110001,
11'b10010110010: edge_mask_reg_512p4[210] <= 1'b1;
 		default: edge_mask_reg_512p4[210] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b1001100010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1101100001,
11'b1101100010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001110001,
11'b10001110010: edge_mask_reg_512p4[211] <= 1'b1;
 		default: edge_mask_reg_512p4[211] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110010,
11'b10110110011,
11'b10110110100: edge_mask_reg_512p4[212] <= 1'b1;
 		default: edge_mask_reg_512p4[212] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001010,
11'b1000110101,
11'b1000110110,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100110011,
11'b10100110100,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100101,
11'b10101100110: edge_mask_reg_512p4[213] <= 1'b1;
 		default: edge_mask_reg_512p4[213] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100111,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000010,
11'b1110000011,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[214] <= 1'b1;
 		default: edge_mask_reg_512p4[214] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000101,
11'b11010000110,
11'b11101010011,
11'b11101100011,
11'b11101100100,
11'b11101110011,
11'b11101110100: edge_mask_reg_512p4[215] <= 1'b1;
 		default: edge_mask_reg_512p4[215] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110000,
11'b10110001,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110010100,
11'b1110010101,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100: edge_mask_reg_512p4[216] <= 1'b1;
 		default: edge_mask_reg_512p4[216] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[217] <= 1'b1;
 		default: edge_mask_reg_512p4[217] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010000,
11'b1101010010,
11'b1101010011,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[218] <= 1'b1;
 		default: edge_mask_reg_512p4[218] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[219] <= 1'b1;
 		default: edge_mask_reg_512p4[219] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110111,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11110000110,
11'b11110010101,
11'b11110010110,
11'b11110100101,
11'b11110100110,
11'b11110110101: edge_mask_reg_512p4[220] <= 1'b1;
 		default: edge_mask_reg_512p4[220] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110001000,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[221] <= 1'b1;
 		default: edge_mask_reg_512p4[221] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000111,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101010001,
11'b1101010010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100001,
11'b1101100010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110110,
11'b1101110111,
11'b1101111000: edge_mask_reg_512p4[222] <= 1'b1;
 		default: edge_mask_reg_512p4[222] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000010,
11'b1111000011: edge_mask_reg_512p4[223] <= 1'b1;
 		default: edge_mask_reg_512p4[223] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100011,
11'b1101100100,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010: edge_mask_reg_512p4[224] <= 1'b1;
 		default: edge_mask_reg_512p4[224] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b101111001,
11'b101111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10110110011,
11'b10110110100,
11'b10111000100: edge_mask_reg_512p4[225] <= 1'b1;
 		default: edge_mask_reg_512p4[225] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000011,
11'b1011000100,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10111000100: edge_mask_reg_512p4[226] <= 1'b1;
 		default: edge_mask_reg_512p4[226] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011010011,
11'b1011010100,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111010011,
11'b1111010100,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10111000100: edge_mask_reg_512p4[227] <= 1'b1;
 		default: edge_mask_reg_512p4[227] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001100011,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011: edge_mask_reg_512p4[228] <= 1'b1;
 		default: edge_mask_reg_512p4[228] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1100010011,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110: edge_mask_reg_512p4[229] <= 1'b1;
 		default: edge_mask_reg_512p4[229] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[230] <= 1'b1;
 		default: edge_mask_reg_512p4[230] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[231] <= 1'b1;
 		default: edge_mask_reg_512p4[231] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b11001010010,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11101010011,
11'b11101010100,
11'b11101010101,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101110100: edge_mask_reg_512p4[232] <= 1'b1;
 		default: edge_mask_reg_512p4[232] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101101000: edge_mask_reg_512p4[233] <= 1'b1;
 		default: edge_mask_reg_512p4[233] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000010,
11'b101000011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101101000: edge_mask_reg_512p4[234] <= 1'b1;
 		default: edge_mask_reg_512p4[234] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011001,
11'b10001100011,
11'b10001100100,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10110000001,
11'b10110010001: edge_mask_reg_512p4[235] <= 1'b1;
 		default: edge_mask_reg_512p4[235] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b1000110100,
11'b1000110101,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100110100,
11'b1100110101,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100011,
11'b10001100100,
11'b10001100101: edge_mask_reg_512p4[236] <= 1'b1;
 		default: edge_mask_reg_512p4[236] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110100,
11'b10010010100,
11'b10010010101,
11'b10010100100,
11'b10010100101: edge_mask_reg_512p4[237] <= 1'b1;
 		default: edge_mask_reg_512p4[237] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[238] <= 1'b1;
 		default: edge_mask_reg_512p4[238] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[239] <= 1'b1;
 		default: edge_mask_reg_512p4[239] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b101011001,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000111,
11'b10010001000,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101100100,
11'b11101110100,
11'b11101110101,
11'b11110000100: edge_mask_reg_512p4[240] <= 1'b1;
 		default: edge_mask_reg_512p4[240] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11101110100,
11'b11110000100: edge_mask_reg_512p4[241] <= 1'b1;
 		default: edge_mask_reg_512p4[241] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100001,
11'b11100010,
11'b11100011,
11'b11100100,
11'b11100101,
11'b110111000,
11'b111000001,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111100011,
11'b111100100: edge_mask_reg_512p4[242] <= 1'b1;
 		default: edge_mask_reg_512p4[242] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100111,
11'b101101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100111,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[243] <= 1'b1;
 		default: edge_mask_reg_512p4[243] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110010,
11'b10110110011,
11'b10110110100: edge_mask_reg_512p4[244] <= 1'b1;
 		default: edge_mask_reg_512p4[244] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[245] <= 1'b1;
 		default: edge_mask_reg_512p4[245] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11110011,
11'b11110100,
11'b11110101: edge_mask_reg_512p4[246] <= 1'b1;
 		default: edge_mask_reg_512p4[246] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111000,
11'b10111001,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100100,
11'b11100101,
11'b11100110: edge_mask_reg_512p4[247] <= 1'b1;
 		default: edge_mask_reg_512p4[247] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1110000010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110000,
11'b10010110001: edge_mask_reg_512p4[248] <= 1'b1;
 		default: edge_mask_reg_512p4[248] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100011,
11'b100100,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100011,
11'b100100100,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100110001,
11'b1100110010,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010011,
11'b1101010100,
11'b1101010101: edge_mask_reg_512p4[249] <= 1'b1;
 		default: edge_mask_reg_512p4[249] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111001,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101: edge_mask_reg_512p4[250] <= 1'b1;
 		default: edge_mask_reg_512p4[250] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11110000100,
11'b11110000101,
11'b11110000110,
11'b11110000111,
11'b11110001000,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110010111,
11'b11110011000: edge_mask_reg_512p4[251] <= 1'b1;
 		default: edge_mask_reg_512p4[251] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110101,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010011,
11'b1101010100,
11'b1101010101: edge_mask_reg_512p4[252] <= 1'b1;
 		default: edge_mask_reg_512p4[252] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010: edge_mask_reg_512p4[253] <= 1'b1;
 		default: edge_mask_reg_512p4[253] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b111000,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000,
11'b1011001: edge_mask_reg_512p4[254] <= 1'b1;
 		default: edge_mask_reg_512p4[254] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10101010001,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101100000,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p4[255] <= 1'b1;
 		default: edge_mask_reg_512p4[255] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000010,
11'b1110010101,
11'b1110010110,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000010: edge_mask_reg_512p4[256] <= 1'b1;
 		default: edge_mask_reg_512p4[256] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011: edge_mask_reg_512p4[257] <= 1'b1;
 		default: edge_mask_reg_512p4[257] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010: edge_mask_reg_512p4[258] <= 1'b1;
 		default: edge_mask_reg_512p4[258] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[259] <= 1'b1;
 		default: edge_mask_reg_512p4[259] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110010,
11'b10001110011,
11'b10101010000,
11'b10101010001,
11'b10101100000,
11'b10101100001: edge_mask_reg_512p4[260] <= 1'b1;
 		default: edge_mask_reg_512p4[260] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100010,
11'b10001100011,
11'b10001100100: edge_mask_reg_512p4[261] <= 1'b1;
 		default: edge_mask_reg_512p4[261] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110011,
11'b10110110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110011,
11'b11110010100: edge_mask_reg_512p4[262] <= 1'b1;
 		default: edge_mask_reg_512p4[262] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110101,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b10000110001,
11'b10001000000,
11'b10001000001,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100: edge_mask_reg_512p4[263] <= 1'b1;
 		default: edge_mask_reg_512p4[263] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101: edge_mask_reg_512p4[264] <= 1'b1;
 		default: edge_mask_reg_512p4[264] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010111000,
11'b1010111001,
11'b1110100011: edge_mask_reg_512p4[265] <= 1'b1;
 		default: edge_mask_reg_512p4[265] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110010,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110110001,
11'b10110110010: edge_mask_reg_512p4[266] <= 1'b1;
 		default: edge_mask_reg_512p4[266] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p4[267] <= 1'b1;
 		default: edge_mask_reg_512p4[267] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b10001100010: edge_mask_reg_512p4[268] <= 1'b1;
 		default: edge_mask_reg_512p4[268] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[269] <= 1'b1;
 		default: edge_mask_reg_512p4[269] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110110001,
11'b10110110010: edge_mask_reg_512p4[270] <= 1'b1;
 		default: edge_mask_reg_512p4[270] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100: edge_mask_reg_512p4[271] <= 1'b1;
 		default: edge_mask_reg_512p4[271] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011,
11'b10110000010,
11'b10110000011,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100: edge_mask_reg_512p4[272] <= 1'b1;
 		default: edge_mask_reg_512p4[272] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000,
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b110100,
11'b110111,
11'b111000,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000: edge_mask_reg_512p4[273] <= 1'b1;
 		default: edge_mask_reg_512p4[273] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b110100,
11'b110111,
11'b111000,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010111,
11'b1011000: edge_mask_reg_512p4[274] <= 1'b1;
 		default: edge_mask_reg_512p4[274] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[275] <= 1'b1;
 		default: edge_mask_reg_512p4[275] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[276] <= 1'b1;
 		default: edge_mask_reg_512p4[276] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[277] <= 1'b1;
 		default: edge_mask_reg_512p4[277] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011: edge_mask_reg_512p4[278] <= 1'b1;
 		default: edge_mask_reg_512p4[278] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000000,
11'b1111000001,
11'b1111000010,
11'b1111000011: edge_mask_reg_512p4[279] <= 1'b1;
 		default: edge_mask_reg_512p4[279] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[280] <= 1'b1;
 		default: edge_mask_reg_512p4[280] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101: edge_mask_reg_512p4[281] <= 1'b1;
 		default: edge_mask_reg_512p4[281] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001000110: edge_mask_reg_512p4[282] <= 1'b1;
 		default: edge_mask_reg_512p4[282] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110010011,
11'b1110010100,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[283] <= 1'b1;
 		default: edge_mask_reg_512p4[283] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[284] <= 1'b1;
 		default: edge_mask_reg_512p4[284] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11101100100,
11'b11101100101,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000011,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[285] <= 1'b1;
 		default: edge_mask_reg_512p4[285] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11011001,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11110100,
11'b11110101,
11'b11110110,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111100111,
11'b111101000,
11'b111110100,
11'b111110101,
11'b111110110,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011110101,
11'b1011110110,
11'b1111010110,
11'b1111010111,
11'b1111100101,
11'b1111100110,
11'b1111110101,
11'b1111110110: edge_mask_reg_512p4[286] <= 1'b1;
 		default: edge_mask_reg_512p4[286] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b1111100,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101010,
11'b1101110100,
11'b1101110101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[287] <= 1'b1;
 		default: edge_mask_reg_512p4[287] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b101011000,
11'b101011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[288] <= 1'b1;
 		default: edge_mask_reg_512p4[288] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000111,
11'b111010000,
11'b111010001,
11'b111010010,
11'b111010011,
11'b1010010111,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110111,
11'b1011000001,
11'b1011000010,
11'b1011000011: edge_mask_reg_512p4[289] <= 1'b1;
 		default: edge_mask_reg_512p4[289] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111001,
11'b1001111010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10100110011,
11'b10100110100: edge_mask_reg_512p4[290] <= 1'b1;
 		default: edge_mask_reg_512p4[290] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100110100,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100101,
11'b10101100110: edge_mask_reg_512p4[291] <= 1'b1;
 		default: edge_mask_reg_512p4[291] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p4[292] <= 1'b1;
 		default: edge_mask_reg_512p4[292] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100101,
11'b10101100100,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100011: edge_mask_reg_512p4[293] <= 1'b1;
 		default: edge_mask_reg_512p4[293] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[294] <= 1'b1;
 		default: edge_mask_reg_512p4[294] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010110,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[295] <= 1'b1;
 		default: edge_mask_reg_512p4[295] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p4[296] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100000,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b110000,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100100000,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1001000010,
11'b1001000011,
11'b1001000100: edge_mask_reg_512p4[297] <= 1'b1;
 		default: edge_mask_reg_512p4[297] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100000,
11'b1100001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101101000: edge_mask_reg_512p4[298] <= 1'b1;
 		default: edge_mask_reg_512p4[298] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100011,
11'b1101100100,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b10010000001,
11'b10010000010: edge_mask_reg_512p4[299] <= 1'b1;
 		default: edge_mask_reg_512p4[299] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11110100,
11'b11110101,
11'b11110110,
11'b11110111,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111100111,
11'b111110100,
11'b111110101,
11'b111110110: edge_mask_reg_512p4[300] <= 1'b1;
 		default: edge_mask_reg_512p4[300] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[301] <= 1'b1;
 		default: edge_mask_reg_512p4[301] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[302] <= 1'b1;
 		default: edge_mask_reg_512p4[302] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b110000001,
11'b110000010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p4[303] <= 1'b1;
 		default: edge_mask_reg_512p4[303] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[304] <= 1'b1;
 		default: edge_mask_reg_512p4[304] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010000101,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010110011,
11'b11010110100: edge_mask_reg_512p4[305] <= 1'b1;
 		default: edge_mask_reg_512p4[305] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100001,
11'b1001100010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[306] <= 1'b1;
 		default: edge_mask_reg_512p4[306] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100001,
11'b1001100010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[307] <= 1'b1;
 		default: edge_mask_reg_512p4[307] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b1001100001,
11'b1001100010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1101100011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[308] <= 1'b1;
 		default: edge_mask_reg_512p4[308] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100001,
11'b1001100010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010111,
11'b1110011000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000: edge_mask_reg_512p4[309] <= 1'b1;
 		default: edge_mask_reg_512p4[309] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000: edge_mask_reg_512p4[310] <= 1'b1;
 		default: edge_mask_reg_512p4[310] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000111,
11'b1001001000,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000: edge_mask_reg_512p4[311] <= 1'b1;
 		default: edge_mask_reg_512p4[311] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11100010,
11'b111010010,
11'b111010011: edge_mask_reg_512p4[312] <= 1'b1;
 		default: edge_mask_reg_512p4[312] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100: edge_mask_reg_512p4[313] <= 1'b1;
 		default: edge_mask_reg_512p4[313] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110011,
11'b11010110100: edge_mask_reg_512p4[314] <= 1'b1;
 		default: edge_mask_reg_512p4[314] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[315] <= 1'b1;
 		default: edge_mask_reg_512p4[315] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p4[316] <= 1'b1;
 		default: edge_mask_reg_512p4[316] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100010,
11'b11001110010: edge_mask_reg_512p4[317] <= 1'b1;
 		default: edge_mask_reg_512p4[317] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b11001100010,
11'b11001110010: edge_mask_reg_512p4[318] <= 1'b1;
 		default: edge_mask_reg_512p4[318] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10101010100,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100: edge_mask_reg_512p4[319] <= 1'b1;
 		default: edge_mask_reg_512p4[319] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[320] <= 1'b1;
 		default: edge_mask_reg_512p4[320] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110010,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000010,
11'b10011000011,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b11010100010,
11'b11010100011,
11'b11010100100,
11'b11010110010,
11'b11010110011: edge_mask_reg_512p4[321] <= 1'b1;
 		default: edge_mask_reg_512p4[321] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110111000,
11'b110111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010100001,
11'b10010100010,
11'b10010110001,
11'b10010110010: edge_mask_reg_512p4[322] <= 1'b1;
 		default: edge_mask_reg_512p4[322] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110111000,
11'b110111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110001,
11'b10010110010: edge_mask_reg_512p4[323] <= 1'b1;
 		default: edge_mask_reg_512p4[323] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110111000,
11'b110111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010100001,
11'b10010100010,
11'b10010110001,
11'b10010110010: edge_mask_reg_512p4[324] <= 1'b1;
 		default: edge_mask_reg_512p4[324] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000001,
11'b10000010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100111,
11'b1110101000: edge_mask_reg_512p4[325] <= 1'b1;
 		default: edge_mask_reg_512p4[325] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101: edge_mask_reg_512p4[326] <= 1'b1;
 		default: edge_mask_reg_512p4[326] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b1111100,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b11010010011,
11'b11010010100: edge_mask_reg_512p4[327] <= 1'b1;
 		default: edge_mask_reg_512p4[327] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b1111100,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010100,
11'b11101110100,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[328] <= 1'b1;
 		default: edge_mask_reg_512p4[328] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[329] <= 1'b1;
 		default: edge_mask_reg_512p4[329] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[330] <= 1'b1;
 		default: edge_mask_reg_512p4[330] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110001000,
11'b1110001001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10101100001,
11'b10101100010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[331] <= 1'b1;
 		default: edge_mask_reg_512p4[331] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10010100110,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100011,
11'b10110100101,
11'b10110100110,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11110000100,
11'b11110010100: edge_mask_reg_512p4[332] <= 1'b1;
 		default: edge_mask_reg_512p4[332] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111000,
11'b10111001,
11'b11010100,
11'b11010101,
11'b11100100,
11'b11100101: edge_mask_reg_512p4[333] <= 1'b1;
 		default: edge_mask_reg_512p4[333] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100010,
11'b100011,
11'b110000,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b101000111,
11'b101001000,
11'b101010111,
11'b101011000: edge_mask_reg_512p4[334] <= 1'b1;
 		default: edge_mask_reg_512p4[334] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100011,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101: edge_mask_reg_512p4[335] <= 1'b1;
 		default: edge_mask_reg_512p4[335] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[336] <= 1'b1;
 		default: edge_mask_reg_512p4[336] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100111,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[337] <= 1'b1;
 		default: edge_mask_reg_512p4[337] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101110001,
11'b10101110010: edge_mask_reg_512p4[338] <= 1'b1;
 		default: edge_mask_reg_512p4[338] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010010011,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p4[339] <= 1'b1;
 		default: edge_mask_reg_512p4[339] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b110000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000: edge_mask_reg_512p4[340] <= 1'b1;
 		default: edge_mask_reg_512p4[340] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b110000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000: edge_mask_reg_512p4[341] <= 1'b1;
 		default: edge_mask_reg_512p4[341] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110000010,
11'b1110000011,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110110010,
11'b1110110011: edge_mask_reg_512p4[342] <= 1'b1;
 		default: edge_mask_reg_512p4[342] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101: edge_mask_reg_512p4[343] <= 1'b1;
 		default: edge_mask_reg_512p4[343] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110010,
11'b10110110011: edge_mask_reg_512p4[344] <= 1'b1;
 		default: edge_mask_reg_512p4[344] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110010000,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100000,
11'b10110100001,
11'b10110100010,
11'b10110100011: edge_mask_reg_512p4[345] <= 1'b1;
 		default: edge_mask_reg_512p4[345] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010011,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000110: edge_mask_reg_512p4[346] <= 1'b1;
 		default: edge_mask_reg_512p4[346] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100110000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000110000,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001001000,
11'b1001001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001111000,
11'b1001111001,
11'b1100110000,
11'b1100110001,
11'b1101000000,
11'b1101000001,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110: edge_mask_reg_512p4[347] <= 1'b1;
 		default: edge_mask_reg_512p4[347] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[348] <= 1'b1;
 		default: edge_mask_reg_512p4[348] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010000,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[349] <= 1'b1;
 		default: edge_mask_reg_512p4[349] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110: edge_mask_reg_512p4[350] <= 1'b1;
 		default: edge_mask_reg_512p4[350] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101010011,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000010,
11'b11010000011,
11'b11010000100: edge_mask_reg_512p4[351] <= 1'b1;
 		default: edge_mask_reg_512p4[351] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001100111,
11'b1001101000,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[352] <= 1'b1;
 		default: edge_mask_reg_512p4[352] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[353] <= 1'b1;
 		default: edge_mask_reg_512p4[353] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b10001110010,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p4[354] <= 1'b1;
 		default: edge_mask_reg_512p4[354] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[355] <= 1'b1;
 		default: edge_mask_reg_512p4[355] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b1110011001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[356] <= 1'b1;
 		default: edge_mask_reg_512p4[356] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b10010000000,
11'b10010000001,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[357] <= 1'b1;
 		default: edge_mask_reg_512p4[357] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101101000,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b10010000000,
11'b10010000001,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[358] <= 1'b1;
 		default: edge_mask_reg_512p4[358] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1011000011: edge_mask_reg_512p4[359] <= 1'b1;
 		default: edge_mask_reg_512p4[359] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000010,
11'b1011000011,
11'b1011000100: edge_mask_reg_512p4[360] <= 1'b1;
 		default: edge_mask_reg_512p4[360] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1111000001,
11'b1111000010: edge_mask_reg_512p4[361] <= 1'b1;
 		default: edge_mask_reg_512p4[361] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b11001100001,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110001,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11010000001,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010010011,
11'b11010010100,
11'b11101100001,
11'b11101110001: edge_mask_reg_512p4[362] <= 1'b1;
 		default: edge_mask_reg_512p4[362] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[363] <= 1'b1;
 		default: edge_mask_reg_512p4[363] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[364] <= 1'b1;
 		default: edge_mask_reg_512p4[364] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[365] <= 1'b1;
 		default: edge_mask_reg_512p4[365] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[366] <= 1'b1;
 		default: edge_mask_reg_512p4[366] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[367] <= 1'b1;
 		default: edge_mask_reg_512p4[367] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100010,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[368] <= 1'b1;
 		default: edge_mask_reg_512p4[368] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100111,
11'b1110101000,
11'b1110101001: edge_mask_reg_512p4[369] <= 1'b1;
 		default: edge_mask_reg_512p4[369] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110111,
11'b1010111000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010: edge_mask_reg_512p4[370] <= 1'b1;
 		default: edge_mask_reg_512p4[370] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010: edge_mask_reg_512p4[371] <= 1'b1;
 		default: edge_mask_reg_512p4[371] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100: edge_mask_reg_512p4[372] <= 1'b1;
 		default: edge_mask_reg_512p4[372] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[373] <= 1'b1;
 		default: edge_mask_reg_512p4[373] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1110010001,
11'b1110010010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010: edge_mask_reg_512p4[374] <= 1'b1;
 		default: edge_mask_reg_512p4[374] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[375] <= 1'b1;
 		default: edge_mask_reg_512p4[375] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1110000111,
11'b1110001000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110000,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[376] <= 1'b1;
 		default: edge_mask_reg_512p4[376] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11100010,
11'b11100011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b111100010,
11'b111100011: edge_mask_reg_512p4[377] <= 1'b1;
 		default: edge_mask_reg_512p4[377] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10010000011,
11'b10010000100,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011: edge_mask_reg_512p4[378] <= 1'b1;
 		default: edge_mask_reg_512p4[378] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101001,
11'b1010101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10110000010,
11'b10110010010: edge_mask_reg_512p4[379] <= 1'b1;
 		default: edge_mask_reg_512p4[379] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110100,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b10001110011,
11'b10001110100,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100: edge_mask_reg_512p4[380] <= 1'b1;
 		default: edge_mask_reg_512p4[380] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[381] <= 1'b1;
 		default: edge_mask_reg_512p4[381] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b1111100,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101010,
11'b10101011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100100,
11'b10110100101,
11'b10110100110: edge_mask_reg_512p4[382] <= 1'b1;
 		default: edge_mask_reg_512p4[382] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110: edge_mask_reg_512p4[383] <= 1'b1;
 		default: edge_mask_reg_512p4[383] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10101010101,
11'b10101010110,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11101110011: edge_mask_reg_512p4[384] <= 1'b1;
 		default: edge_mask_reg_512p4[384] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101110011: edge_mask_reg_512p4[385] <= 1'b1;
 		default: edge_mask_reg_512p4[385] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000101,
11'b11101010100,
11'b11101010101,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101110011,
11'b11101110100: edge_mask_reg_512p4[386] <= 1'b1;
 		default: edge_mask_reg_512p4[386] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101100001,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11010000010: edge_mask_reg_512p4[387] <= 1'b1;
 		default: edge_mask_reg_512p4[387] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100010001,
11'b100010010,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010001,
11'b1000010010,
11'b1000010011,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001011000,
11'b1001011001,
11'b1001101000,
11'b1001101001,
11'b1100010010,
11'b1100010011,
11'b1100100010,
11'b1100100011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b10000100011: edge_mask_reg_512p4[388] <= 1'b1;
 		default: edge_mask_reg_512p4[388] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000,
11'b10010010001: edge_mask_reg_512p4[389] <= 1'b1;
 		default: edge_mask_reg_512p4[389] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11011001,
11'b11011010,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11101001,
11'b11110100,
11'b11110101,
11'b11110110,
11'b11110111,
11'b11111000,
11'b110101001,
11'b110101010,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111100101,
11'b111100110,
11'b111100111,
11'b111101000,
11'b111101001,
11'b111110101,
11'b111110110,
11'b111110111,
11'b111111000,
11'b1011001000,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011110110,
11'b1011110111,
11'b1011111000: edge_mask_reg_512p4[390] <= 1'b1;
 		default: edge_mask_reg_512p4[390] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11,
11'b100,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b10111,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100010101,
11'b100010110,
11'b100100101,
11'b100100110: edge_mask_reg_512p4[391] <= 1'b1;
 		default: edge_mask_reg_512p4[391] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[392] <= 1'b1;
 		default: edge_mask_reg_512p4[392] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[393] <= 1'b1;
 		default: edge_mask_reg_512p4[393] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[394] <= 1'b1;
 		default: edge_mask_reg_512p4[394] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[395] <= 1'b1;
 		default: edge_mask_reg_512p4[395] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[396] <= 1'b1;
 		default: edge_mask_reg_512p4[396] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[397] <= 1'b1;
 		default: edge_mask_reg_512p4[397] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101010101,
11'b101010110,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010011,
11'b1101010100,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000001,
11'b1110000010,
11'b1110001000,
11'b1110001001,
11'b10001100001,
11'b10001100010,
11'b10001110001,
11'b10001110010: edge_mask_reg_512p4[398] <= 1'b1;
 		default: edge_mask_reg_512p4[398] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110100,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[399] <= 1'b1;
 		default: edge_mask_reg_512p4[399] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10010000010,
11'b10010010010: edge_mask_reg_512p4[400] <= 1'b1;
 		default: edge_mask_reg_512p4[400] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[401] <= 1'b1;
 		default: edge_mask_reg_512p4[401] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1110001000,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110001,
11'b10010110010,
11'b10010110011: edge_mask_reg_512p4[402] <= 1'b1;
 		default: edge_mask_reg_512p4[402] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b1010000111,
11'b1010001000,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1110010010,
11'b1110010011,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110110010,
11'b1110110011: edge_mask_reg_512p4[403] <= 1'b1;
 		default: edge_mask_reg_512p4[403] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010: edge_mask_reg_512p4[404] <= 1'b1;
 		default: edge_mask_reg_512p4[404] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[405] <= 1'b1;
 		default: edge_mask_reg_512p4[405] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[406] <= 1'b1;
 		default: edge_mask_reg_512p4[406] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[407] <= 1'b1;
 		default: edge_mask_reg_512p4[407] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100010,
11'b1100011,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110010,
11'b1110011,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[408] <= 1'b1;
 		default: edge_mask_reg_512p4[408] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[409] <= 1'b1;
 		default: edge_mask_reg_512p4[409] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001: edge_mask_reg_512p4[410] <= 1'b1;
 		default: edge_mask_reg_512p4[410] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[411] <= 1'b1;
 		default: edge_mask_reg_512p4[411] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11001000,
11'b11010011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[412] <= 1'b1;
 		default: edge_mask_reg_512p4[412] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[413] <= 1'b1;
 		default: edge_mask_reg_512p4[413] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[414] <= 1'b1;
 		default: edge_mask_reg_512p4[414] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010001,
11'b111010010,
11'b111010011,
11'b111010100,
11'b111010101,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011010001,
11'b1011010010,
11'b1011010011,
11'b1011010100,
11'b1011010101,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011,
11'b1111000100: edge_mask_reg_512p4[415] <= 1'b1;
 		default: edge_mask_reg_512p4[415] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[416] <= 1'b1;
 		default: edge_mask_reg_512p4[416] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b10001110011,
11'b10001110100,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[417] <= 1'b1;
 		default: edge_mask_reg_512p4[417] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011: edge_mask_reg_512p4[418] <= 1'b1;
 		default: edge_mask_reg_512p4[418] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001000010,
11'b1001000011,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b10001010000,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011: edge_mask_reg_512p4[419] <= 1'b1;
 		default: edge_mask_reg_512p4[419] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101001000,
11'b101001001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001000010,
11'b1001000011,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b10001010000,
11'b10001010001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011: edge_mask_reg_512p4[420] <= 1'b1;
 		default: edge_mask_reg_512p4[420] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101001000,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001000010,
11'b1001000011,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000010,
11'b1101000011,
11'b1101010000,
11'b1101010001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b10001010000,
11'b10001010001,
11'b10001010010,
11'b10001010011,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011: edge_mask_reg_512p4[421] <= 1'b1;
 		default: edge_mask_reg_512p4[421] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011: edge_mask_reg_512p4[422] <= 1'b1;
 		default: edge_mask_reg_512p4[422] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100: edge_mask_reg_512p4[423] <= 1'b1;
 		default: edge_mask_reg_512p4[423] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11110000100,
11'b11110010100: edge_mask_reg_512p4[424] <= 1'b1;
 		default: edge_mask_reg_512p4[424] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[425] <= 1'b1;
 		default: edge_mask_reg_512p4[425] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b11001010110,
11'b11001010111,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000011,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p4[426] <= 1'b1;
 		default: edge_mask_reg_512p4[426] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1101100001,
11'b1101100010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[427] <= 1'b1;
 		default: edge_mask_reg_512p4[427] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1101100001,
11'b1101100010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000001,
11'b1110000010,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[428] <= 1'b1;
 		default: edge_mask_reg_512p4[428] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100100,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001: edge_mask_reg_512p4[429] <= 1'b1;
 		default: edge_mask_reg_512p4[429] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110010,
11'b110111,
11'b111000,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010100,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b100110000,
11'b101000000,
11'b101000001,
11'b101000010,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1001000000,
11'b1001000001,
11'b1001000010,
11'b1001000011,
11'b1001000100,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000: edge_mask_reg_512p4[430] <= 1'b1;
 		default: edge_mask_reg_512p4[430] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100010,
11'b100011,
11'b110000,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000000,
11'b1000001,
11'b1000010,
11'b1000011,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b100110001,
11'b100110010,
11'b100110011,
11'b101000111,
11'b101001000,
11'b101010111,
11'b101011000: edge_mask_reg_512p4[431] <= 1'b1;
 		default: edge_mask_reg_512p4[431] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p4[432] <= 1'b1;
 		default: edge_mask_reg_512p4[432] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001: edge_mask_reg_512p4[433] <= 1'b1;
 		default: edge_mask_reg_512p4[433] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b10001100001,
11'b10001100010,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10010000000: edge_mask_reg_512p4[434] <= 1'b1;
 		default: edge_mask_reg_512p4[434] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011001,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p4[435] <= 1'b1;
 		default: edge_mask_reg_512p4[435] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110111,
11'b1010111000: edge_mask_reg_512p4[436] <= 1'b1;
 		default: edge_mask_reg_512p4[436] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1110010101,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110: edge_mask_reg_512p4[437] <= 1'b1;
 		default: edge_mask_reg_512p4[437] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110100,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110100,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101: edge_mask_reg_512p4[438] <= 1'b1;
 		default: edge_mask_reg_512p4[438] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111001,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110001,
11'b10010110100: edge_mask_reg_512p4[439] <= 1'b1;
 		default: edge_mask_reg_512p4[439] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000010,
11'b10000011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010010,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001101000,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[440] <= 1'b1;
 		default: edge_mask_reg_512p4[440] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[441] <= 1'b1;
 		default: edge_mask_reg_512p4[441] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111: edge_mask_reg_512p4[442] <= 1'b1;
 		default: edge_mask_reg_512p4[442] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001001,
11'b1010001010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100110,
11'b11001100111: edge_mask_reg_512p4[443] <= 1'b1;
 		default: edge_mask_reg_512p4[443] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001001,
11'b1010001010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11001100111: edge_mask_reg_512p4[444] <= 1'b1;
 		default: edge_mask_reg_512p4[444] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001001,
11'b1001000110,
11'b1001000111,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10100110101,
11'b10100110110,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b11001000011,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100110: edge_mask_reg_512p4[445] <= 1'b1;
 		default: edge_mask_reg_512p4[445] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10101110001: edge_mask_reg_512p4[446] <= 1'b1;
 		default: edge_mask_reg_512p4[446] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[447] <= 1'b1;
 		default: edge_mask_reg_512p4[447] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100000,
11'b10001100001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000001,
11'b10010000010,
11'b10101110001,
11'b10101110010,
11'b10110000001: edge_mask_reg_512p4[448] <= 1'b1;
 		default: edge_mask_reg_512p4[448] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101110001,
11'b10101110010,
11'b10110000001,
11'b10110000010: edge_mask_reg_512p4[449] <= 1'b1;
 		default: edge_mask_reg_512p4[449] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101110001,
11'b10101110010,
11'b10110000001,
11'b10110000010: edge_mask_reg_512p4[450] <= 1'b1;
 		default: edge_mask_reg_512p4[450] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010111,
11'b10011000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100001,
11'b1001100010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b10001110010,
11'b10001110011,
11'b10010000010: edge_mask_reg_512p4[451] <= 1'b1;
 		default: edge_mask_reg_512p4[451] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p4[452] <= 1'b1;
 		default: edge_mask_reg_512p4[452] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101101000,
11'b1101101001,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10101110001,
11'b10101110011,
11'b10101110100,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101: edge_mask_reg_512p4[453] <= 1'b1;
 		default: edge_mask_reg_512p4[453] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010011,
11'b110010100,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1011000001,
11'b1011000010: edge_mask_reg_512p4[454] <= 1'b1;
 		default: edge_mask_reg_512p4[454] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1011000001,
11'b1011000010,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[455] <= 1'b1;
 		default: edge_mask_reg_512p4[455] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1011000001,
11'b1011000010,
11'b1110010001,
11'b1110010010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100001,
11'b1110100010: edge_mask_reg_512p4[456] <= 1'b1;
 		default: edge_mask_reg_512p4[456] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001,
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110001,
11'b110010,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[457] <= 1'b1;
 		default: edge_mask_reg_512p4[457] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[458] <= 1'b1;
 		default: edge_mask_reg_512p4[458] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100001,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b111010,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[459] <= 1'b1;
 		default: edge_mask_reg_512p4[459] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[460] <= 1'b1;
 		default: edge_mask_reg_512p4[460] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100010,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100010010,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[461] <= 1'b1;
 		default: edge_mask_reg_512p4[461] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11,
11'b100,
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100000011,
11'b100000100,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010011,
11'b1000010100,
11'b1000100101,
11'b1000100110: edge_mask_reg_512p4[462] <= 1'b1;
 		default: edge_mask_reg_512p4[462] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000100,
11'b11110000101,
11'b11110000110,
11'b11110010100,
11'b11110010101: edge_mask_reg_512p4[463] <= 1'b1;
 		default: edge_mask_reg_512p4[463] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100001,
11'b1110100010,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100001,
11'b10010100010,
11'b10110000011,
11'b10110000100,
11'b10110010001,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110100001,
11'b10110100010: edge_mask_reg_512p4[464] <= 1'b1;
 		default: edge_mask_reg_512p4[464] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011001000,
11'b1011001001,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110: edge_mask_reg_512p4[465] <= 1'b1;
 		default: edge_mask_reg_512p4[465] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000011,
11'b111000100,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000011,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110110011,
11'b1110110100: edge_mask_reg_512p4[466] <= 1'b1;
 		default: edge_mask_reg_512p4[466] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000011,
11'b111000100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1011000011,
11'b1011000100,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[467] <= 1'b1;
 		default: edge_mask_reg_512p4[467] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[468] <= 1'b1;
 		default: edge_mask_reg_512p4[468] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010110,
11'b1101010111,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11110000100: edge_mask_reg_512p4[469] <= 1'b1;
 		default: edge_mask_reg_512p4[469] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000000,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[470] <= 1'b1;
 		default: edge_mask_reg_512p4[470] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110010,
11'b10010110011,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100001,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110010,
11'b10110110011,
11'b11010010100,
11'b11010100010,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p4[471] <= 1'b1;
 		default: edge_mask_reg_512p4[471] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100010,
11'b100011,
11'b110010,
11'b110011,
11'b110111,
11'b111000,
11'b1000111,
11'b1001000,
11'b1010111,
11'b1011000: edge_mask_reg_512p4[472] <= 1'b1;
 		default: edge_mask_reg_512p4[472] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110011000,
11'b1110011001: edge_mask_reg_512p4[473] <= 1'b1;
 		default: edge_mask_reg_512p4[473] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010000,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b110000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010: edge_mask_reg_512p4[474] <= 1'b1;
 		default: edge_mask_reg_512p4[474] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110001,
11'b10110010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010101000,
11'b1010101001,
11'b1010101010: edge_mask_reg_512p4[475] <= 1'b1;
 		default: edge_mask_reg_512p4[475] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000010,
11'b11000011,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b1010000111,
11'b1010001000,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1110010010,
11'b1110010011,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1111000000,
11'b1111000001: edge_mask_reg_512p4[476] <= 1'b1;
 		default: edge_mask_reg_512p4[476] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p4[477] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1101010110,
11'b1101010111,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[478] <= 1'b1;
 		default: edge_mask_reg_512p4[478] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011,
11'b10100,
11'b10101,
11'b10110,
11'b10111,
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b100111,
11'b101000,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1001011,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b100010011,
11'b100010100,
11'b100010101,
11'b100010110,
11'b100010111,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101001,
11'b101101010,
11'b1000010011,
11'b1000010100,
11'b1000010101,
11'b1000010110,
11'b1000010111,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000111,
11'b1100010100,
11'b1100010101,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100110110,
11'b1100110111: edge_mask_reg_512p4[479] <= 1'b1;
 		default: edge_mask_reg_512p4[479] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010000,
11'b1010001,
11'b1010010,
11'b1010011,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100000,
11'b1100001,
11'b1100010,
11'b1100011,
11'b1100100,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110000,
11'b1110001,
11'b1110010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110110,
11'b1101110111,
11'b1101111000: edge_mask_reg_512p4[480] <= 1'b1;
 		default: edge_mask_reg_512p4[480] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b1001101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[481] <= 1'b1;
 		default: edge_mask_reg_512p4[481] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000001,
11'b10000010,
11'b10000011,
11'b10000100,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010001,
11'b10010010,
11'b10010011,
11'b10010100,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110010,
11'b101110011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001: edge_mask_reg_512p4[482] <= 1'b1;
 		default: edge_mask_reg_512p4[482] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000110101,
11'b1000110110,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000010,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010010,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100110011,
11'b10101000010,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100101,
11'b10101100110: edge_mask_reg_512p4[483] <= 1'b1;
 		default: edge_mask_reg_512p4[483] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b101010000,
11'b101010001,
11'b101010010,
11'b101010011,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100000,
11'b101100001,
11'b101100010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b1001010000,
11'b1001010001,
11'b1001010010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100000,
11'b1001100001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1101010110,
11'b1101010111,
11'b1101100000,
11'b1101100001,
11'b1101100010,
11'b1101100011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000: edge_mask_reg_512p4[484] <= 1'b1;
 		default: edge_mask_reg_512p4[484] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101100111,
11'b1101101000,
11'b1101110000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10001110000,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011: edge_mask_reg_512p4[485] <= 1'b1;
 		default: edge_mask_reg_512p4[485] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10101000101,
11'b10101000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100100,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p4[486] <= 1'b1;
 		default: edge_mask_reg_512p4[486] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10001000101,
11'b10001000110,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10101000101,
11'b10101000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b11001010011,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100100,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p4[487] <= 1'b1;
 		default: edge_mask_reg_512p4[487] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000110,
11'b10010000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110011,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100011,
11'b11101100100,
11'b11101100101,
11'b11101100110,
11'b11101110011,
11'b11101110100,
11'b11101110101,
11'b11110000100: edge_mask_reg_512p4[488] <= 1'b1;
 		default: edge_mask_reg_512p4[488] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10001100,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10011100,
11'b10101001,
11'b10101010,
11'b10101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110: edge_mask_reg_512p4[489] <= 1'b1;
 		default: edge_mask_reg_512p4[489] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101,
11'b110100111,
11'b110110111,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111010001,
11'b111010010,
11'b111010011: edge_mask_reg_512p4[490] <= 1'b1;
 		default: edge_mask_reg_512p4[490] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000000,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000101,
11'b11000111,
11'b11001000,
11'b11010000,
11'b11010001,
11'b11010010,
11'b11010011,
11'b11010100,
11'b11010101: edge_mask_reg_512p4[491] <= 1'b1;
 		default: edge_mask_reg_512p4[491] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[492] <= 1'b1;
 		default: edge_mask_reg_512p4[492] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000: edge_mask_reg_512p4[493] <= 1'b1;
 		default: edge_mask_reg_512p4[493] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101110001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10010000000,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010010000: edge_mask_reg_512p4[494] <= 1'b1;
 		default: edge_mask_reg_512p4[494] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100111,
11'b1101101000,
11'b10000100100,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101: edge_mask_reg_512p4[495] <= 1'b1;
 		default: edge_mask_reg_512p4[495] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000010,
11'b111000011,
11'b1010000111,
11'b1010001000,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1111000001: edge_mask_reg_512p4[496] <= 1'b1;
 		default: edge_mask_reg_512p4[496] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000010,
11'b11000011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000000,
11'b111000001,
11'b111000010,
11'b111000011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000000,
11'b1011000001,
11'b1011000010,
11'b1110100010,
11'b1110100011,
11'b1110110000,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1111000000,
11'b1111000001,
11'b1111000010: edge_mask_reg_512p4[497] <= 1'b1;
 		default: edge_mask_reg_512p4[497] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000101,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11010100,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11110011,
11'b11110100,
11'b11110101,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111010100,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111100011,
11'b111100100,
11'b111100101,
11'b111100110,
11'b111110011,
11'b111110100,
11'b1011010101,
11'b1011010110: edge_mask_reg_512p4[498] <= 1'b1;
 		default: edge_mask_reg_512p4[498] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000110,
11'b10101010010,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000010,
11'b10110000011,
11'b11001100010,
11'b11001100011,
11'b11001100100,
11'b11001100101,
11'b11001110010,
11'b11001110011,
11'b11001110100,
11'b11001110101: edge_mask_reg_512p4[499] <= 1'b1;
 		default: edge_mask_reg_512p4[499] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11110000100,
11'b11110000101,
11'b11110000110,
11'b11110000111,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110010111: edge_mask_reg_512p4[500] <= 1'b1;
 		default: edge_mask_reg_512p4[500] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1011000001,
11'b1011000010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110110001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1111000001,
11'b1111000010,
11'b1111000011: edge_mask_reg_512p4[501] <= 1'b1;
 		default: edge_mask_reg_512p4[501] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100011,
11'b100100,
11'b100101,
11'b100110,
11'b110011,
11'b110100,
11'b110101,
11'b110110,
11'b110111,
11'b111000,
11'b111001,
11'b1000100,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100010001,
11'b100010010,
11'b100100001,
11'b100100010,
11'b100100011,
11'b100100100,
11'b100100101,
11'b100100110,
11'b100110001,
11'b100110010,
11'b100110011,
11'b100110100,
11'b100110101,
11'b100110110,
11'b100110111,
11'b101000011,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010001,
11'b1000010010,
11'b1000100001,
11'b1000100010,
11'b1000100011,
11'b1000100100,
11'b1000100101,
11'b1000110001,
11'b1000110010,
11'b1000110011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001101000,
11'b1001101001,
11'b1100100001,
11'b1100100010,
11'b1100100011,
11'b1100110001,
11'b1100110010,
11'b1100110011,
11'b1100110100,
11'b1101000011,
11'b1101000100,
11'b1101000101: edge_mask_reg_512p4[502] <= 1'b1;
 		default: edge_mask_reg_512p4[502] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11010101,
11'b11010110,
11'b11010111,
11'b11011000,
11'b11100011,
11'b11100100,
11'b11100101,
11'b11100110,
11'b11100111,
11'b11101000,
11'b11110011,
11'b11110100,
11'b11110101,
11'b11110110,
11'b11110111: edge_mask_reg_512p4[503] <= 1'b1;
 		default: edge_mask_reg_512p4[503] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101000,
11'b10101001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010010,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100010,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11010000010,
11'b11010000011,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010010,
11'b11010010011,
11'b11010010100,
11'b11010010101,
11'b11010100010,
11'b11010100011,
11'b11010100100: edge_mask_reg_512p4[504] <= 1'b1;
 		default: edge_mask_reg_512p4[504] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010011,
11'b110010100,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000111,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1011000010: edge_mask_reg_512p4[505] <= 1'b1;
 		default: edge_mask_reg_512p4[505] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100000,
11'b10100001,
11'b10100010,
11'b10100011,
11'b10100100,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110000,
11'b10110001,
11'b10110010,
11'b10110011,
11'b10110100,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000001,
11'b11000010,
11'b11000011,
11'b11000100,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100001,
11'b110100010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110000,
11'b110110001,
11'b110110010,
11'b110110011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000001,
11'b111000010,
11'b111000011,
11'b111000100,
11'b111000111,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110000,
11'b1010110001,
11'b1010110010,
11'b1010110011,
11'b1010110100,
11'b1010110111,
11'b1010111000,
11'b1011000001,
11'b1011000010: edge_mask_reg_512p4[506] <= 1'b1;
 		default: edge_mask_reg_512p4[506] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b101110001,
11'b101110010,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p4[507] <= 1'b1;
 		default: edge_mask_reg_512p4[507] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1110000010,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110110000,
11'b1110110001,
11'b10010010000,
11'b10010010001,
11'b10010010010,
11'b10010010011,
11'b10010010100,
11'b10010100000,
11'b10010100001,
11'b10010100010,
11'b10010100011,
11'b10010100100: edge_mask_reg_512p4[508] <= 1'b1;
 		default: edge_mask_reg_512p4[508] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b101110011,
11'b101110100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000000,
11'b110000001,
11'b110000010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010000,
11'b110010001,
11'b110010010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001110001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000000,
11'b1010000001,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010000,
11'b1010010001,
11'b1010010010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100000,
11'b1010100001,
11'b1010100010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000000,
11'b1110000001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010000,
11'b1110010001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100000,
11'b1110100001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b10010000001,
11'b10010000010,
11'b10010010001,
11'b10010010010: edge_mask_reg_512p4[509] <= 1'b1;
 		default: edge_mask_reg_512p4[509] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b101011000,
11'b101011001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b1001011000,
11'b1001011001,
11'b1001100010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b10001100010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110001,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000001,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10101100010,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b11001110010,
11'b11010000010: edge_mask_reg_512p4[510] <= 1'b1;
 		default: edge_mask_reg_512p4[510] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110010,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010010,
11'b10010010011,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110001,
11'b10101110010,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000001,
11'b10110000010,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010010,
11'b10110010011,
11'b11001110010,
11'b11001110011,
11'b11010000010,
11'b11010000011: edge_mask_reg_512p4[511] <= 1'b1;
 		default: edge_mask_reg_512p4[511] <= 1'b0;
 	endcase

end
endmodule

